// ------------------------------------------------------------
// Company           :   racyics                      
// Author            :   schreiter            
// E-Mail            :   schreiter@racyics.com                    
//                                      
// Filename          :                   
// Project Name      :   p_ri
// Subproject Name   :   s_libio_gf22fdsoi
// Description       :               
//
// Create Date       :   Wed Sep 12 16:32:15 2018 
// Last Change       :   $Date: 2020-08-20 10:35:38 +0200 (Thu, 20 Aug 2020) $
// by                :   $Author: henker $                                      
// ------------------------------------------------------------
`celldefine
module RIIO_BOND60_INNER_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60_INNER_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60_INNER_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60_OUTER_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60_OUTER_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60_OUTER_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60_PLAIN_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60_PLAIN_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60_PLAIN_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_INNER_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_INNER_GND_CESD( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_INNER_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_INNER_PWR_CESD( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_INNER_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_INNER_SIG_CESD( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_OUTER_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_OUTER_GND_CESD( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_OUTER_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_OUTER_PWR_CESD( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_OUTER_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_OUTER_SIG_CESD( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_PLAIN_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_PLAIN_GND_CESD( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_PLAIN_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_PLAIN_PWR_CESD( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_PLAIN_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND60x90_PLAIN_SIG_CESD( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND64_INNER_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND64_INNER_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND64_INNER_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND64_OUTER_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND64_OUTER_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND64_OUTER_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND64_PLAIN_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND64_PLAIN_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND64_PLAIN_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND70_INNER_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND70_INNER_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND70_INNER_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND70_OUTER_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND70_OUTER_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND70_OUTER_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND70_PLAIN_GND( VSS);
    inout VSS;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND70_PLAIN_PWR( VDD);
    inout VDD;
endmodule
`endcelldefine
`celldefine
module RIIO_BOND70_PLAIN_SIG( PAD);
    inout PAD;
endmodule
`endcelldefine
