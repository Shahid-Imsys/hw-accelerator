-- NoC register Part of NoC simulation pkg
-- 
-- Design: Harald bergh
-- Implemented: Bengt Andersson
-- Revision 0

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library work;
use work.defines.all;

entity NoC_ctrl is
port (
		
		NoCbus	: out std_logic_vector (511 downto 0);
	
);
end NoC_ctrl;


architecture struct of NoC_ctrl is

begin





end struct NoC_ctrl;