-- IO block simulation for Imsys Accelerator
-- 
-- Top file
-- Design: Imsys AB
-- Implemented: Bengt Andersson
-- Revision 0


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library work;
use work.defines.all;


entity IO_block is
	port (
	);
end IO_block;



architecture struct of IO_block is

end struct IO_block;