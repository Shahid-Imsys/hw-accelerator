VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RIIO_CONN_LB05_GND
  CLASS COVER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_CONN_LB05_GND 0 0 ;
  SIZE 0.5 BY 0.5 ;
  SYMMETRY X Y R90 ;
  PIN SIG
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.204 LAYER LB ;
    PORT
      LAYER LB ;
        RECT 0 0 0.1 0.5 ;
    END
  END SIG
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0.4 0 0.5 0.5 ;
    END
  END VSS
  OBS
    LAYER LB ;
      RECT 0.15 -0.01 0.35 0.51 ;
      RECT 0 0 0.5 0.5 ;
  END
END RIIO_CONN_LB05_GND

MACRO RIIO_CONN_LB05_PWR
  CLASS COVER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_CONN_LB05_PWR 0 0 ;
  SIZE 0.5 BY 0.5 ;
  SYMMETRY X Y R90 ;
  PIN SIG
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.204 LAYER LB ;
    PORT
      LAYER LB ;
        RECT 0 0 0.1 0.5 ;
    END
  END SIG
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0.4 0 0.5 0.5 ;
    END
  END VDD
  OBS
    LAYER LB ;
      RECT 0.15 -0.01 0.35 0.51 ;
      RECT 0 0 0.5 0.5 ;
  END
END RIIO_CONN_LB05_PWR

MACRO RIIO_EG1D80V_ESD_B2B_010x046
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ESD_B2B_010x046 0 0 ;
  SIZE 10 BY 46 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER C1 ;
        RECT 0.25 0 0.75 46 ;
    END
    PORT
      LAYER C1 ;
        RECT 1.75 0 2.25 46 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.25 0 3.75 46 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.25 0 6.75 46 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.75 0 8.25 46 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.25 0 9.75 46 ;
    END
  END VSS
  PIN SUB
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "sub SUB!" ;
    PORT
      LAYER C1 ;
        RECT 4.75 0 5.25 46 ;
    END
  END SUB
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER C1 ;
        RECT 1 0.125 1.5 45.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.5 0.125 3 45.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 4 0.125 4.5 45.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.5 0.125 6 45.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 7 0.125 7.5 45.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.5 0.125 9 45.875 ;
    END
  END VSSX
  OBS
    LAYER CA ;
      RECT 0 0 10 46 ;
    LAYER M1 ;
      RECT 0 0 10 46 ;
    LAYER V1 ;
      RECT 0 0 10 46 ;
    LAYER M2 ;
      RECT 0 0 10 46 ;
    LAYER CB ;
      RECT 0 0 10 46 ;
    LAYER AY ;
      RECT 0 0 10 46 ;
    LAYER C1 ;
      RECT 9.25 0 9.75 46 ;
      RECT 8.5 0.125 9 45.875 ;
      RECT 7.75 0 8.25 46 ;
      RECT 7 0.125 7.5 45.875 ;
      RECT 6.25 0 6.75 46 ;
      RECT 5.5 0.125 6 45.875 ;
      RECT 4.75 0 5.25 46 ;
      RECT 4 0.125 4.5 45.875 ;
      RECT 3.25 0 3.75 46 ;
      RECT 2.5 0.125 3 45.875 ;
      RECT 1.75 0 2.25 46 ;
      RECT 1 0.125 1.5 45.875 ;
      RECT 0.25 0 0.75 46 ;
  END
END RIIO_EG1D80V_ESD_B2B_010x046

MACRO RIIO_EG1D80V_ESD_B2B_012x057
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ESD_B2B_012x057 0 0 ;
  SIZE 12 BY 57.28 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER C1 ;
        RECT 1.625 0 2.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.125 0 3.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 4.625 0 5.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.125 0 6.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.625 0 8.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.125 0 9.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 10.625 0 11.125 57.28 ;
    END
  END VSS
  PIN SUB
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "sub SUB!" ;
    PORT
      LAYER C1 ;
        RECT 0.125 0 0.625 57.28 ;
    END
  END SUB
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER C1 ;
        RECT 0.875 0.125 1.375 57.155 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.375 0.125 2.875 57.155 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.875 0.125 4.375 57.155 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.375 0.125 5.875 57.155 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.875 0.125 7.375 57.155 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.375 0.125 8.875 57.155 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.875 0.125 10.375 57.155 ;
    END
    PORT
      LAYER C1 ;
        RECT 11.375 0.125 11.875 57.155 ;
    END
  END VSSX
  OBS
    LAYER CA ;
      RECT 0 0 12 57.28 ;
    LAYER M1 ;
      RECT 0 0 12 57.28 ;
    LAYER V1 ;
      RECT 0 0 12 57.28 ;
    LAYER M2 ;
      RECT 0 0 12 57.28 ;
    LAYER CB ;
      RECT 0 0 12 57.28 ;
    LAYER AY ;
      RECT 0 0 12 57.28 ;
    LAYER C1 ;
      RECT 11.375 0.125 11.875 57.155 ;
      RECT 10.625 0 11.125 57.28 ;
      RECT 9.875 0.125 10.375 57.155 ;
      RECT 9.125 0 9.625 57.28 ;
      RECT 8.375 0.125 8.875 57.155 ;
      RECT 7.625 0 8.125 57.28 ;
      RECT 6.875 0.125 7.375 57.155 ;
      RECT 6.125 0 6.625 57.28 ;
      RECT 5.375 0.125 5.875 57.155 ;
      RECT 4.625 0 5.125 57.28 ;
      RECT 3.875 0.125 4.375 57.155 ;
      RECT 3.125 0 3.625 57.28 ;
      RECT 2.375 0.125 2.875 57.155 ;
      RECT 1.625 0 2.125 57.28 ;
      RECT 0.875 0.125 1.375 57.155 ;
      RECT 0.125 0 0.625 57.28 ;
  END
END RIIO_EG1D80V_ESD_B2B_012x057

MACRO RIIO_EG1D80V_ESD_B2B_059x010
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ESD_B2B_059x010 0 0 ;
  SIZE 59.25 BY 10 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER C1 ;
        RECT 0.875 0 1.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.375 0 2.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.875 0 4.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.375 0 5.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.875 0 7.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.375 0 8.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.875 0 10.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 11.375 0 11.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 12.875 0 13.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 14.375 0 14.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 15.875 0 16.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 17.375 0 17.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 18.875 0 19.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 20.375 0 20.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 21.875 0 22.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 23.375 0 23.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 24.875 0 25.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 26.375 0 26.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 27.875 0 28.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 29.375 0 29.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 30.875 0 31.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 32.375 0 32.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 33.875 0 34.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 35.375 0 35.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 36.875 0 37.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 38.375 0 38.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 39.875 0 40.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 41.375 0 41.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 42.875 0 43.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 44.375 0 44.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 45.875 0 46.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 47.375 0 47.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 48.875 0 49.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 50.375 0 50.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 51.875 0 52.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 53.375 0 53.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 54.875 0 55.375 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 56.375 0 56.875 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 57.875 0 58.375 10 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER C1 ;
        RECT 1.625 0.125 2.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.125 0.125 3.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 4.625 0.125 5.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.125 0.125 6.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.625 0.125 8.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.125 0.125 9.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 10.625 0.125 11.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 12.125 0.125 12.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 13.625 0.125 14.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 15.125 0.125 15.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 16.625 0.125 17.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 18.125 0.125 18.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 19.625 0.125 20.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 21.125 0.125 21.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 22.625 0.125 23.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 24.125 0.125 24.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 25.625 0.125 26.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 27.125 0.125 27.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 28.625 0.125 29.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 30.125 0.125 30.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 31.625 0.125 32.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 33.125 0.125 33.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 34.625 0.125 35.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 36.125 0.125 36.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 37.625 0.125 38.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 39.125 0.125 39.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 40.625 0.125 41.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 42.125 0.125 42.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 43.625 0.125 44.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 45.125 0.125 45.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 46.625 0.125 47.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 48.125 0.125 48.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 49.625 0.125 50.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 51.125 0.125 51.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 52.625 0.125 53.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 54.125 0.125 54.625 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 55.625 0.125 56.125 9.875 ;
    END
    PORT
      LAYER C1 ;
        RECT 57.125 0.125 57.625 9.875 ;
    END
  END VSSX
  PIN SUB
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "sub SUB!" ;
    PORT
      LAYER C1 ;
        RECT 0.125 0 0.625 10 ;
    END
    PORT
      LAYER C1 ;
        RECT 58.625 0 59.125 10 ;
    END
  END SUB
  OBS
    LAYER CA ;
      RECT 0 0 59.25 10 ;
    LAYER M1 ;
      RECT 0 0 59.25 10 ;
    LAYER V1 ;
      RECT 0 0 59.25 10 ;
    LAYER M2 ;
      RECT 0 0 59.25 10 ;
    LAYER CB ;
      RECT 0 0 59.25 10 ;
    LAYER AY ;
      RECT 0 0 59.25 10 ;
    LAYER C1 ;
      RECT 58.625 0 59.125 10 ;
      RECT 57.875 0 58.375 10 ;
      RECT 57.125 0.125 57.625 9.875 ;
      RECT 56.375 0 56.875 10 ;
      RECT 55.625 0.125 56.125 9.875 ;
      RECT 54.875 0 55.375 10 ;
      RECT 54.125 0.125 54.625 9.875 ;
      RECT 53.375 0 53.875 10 ;
      RECT 52.625 0.125 53.125 9.875 ;
      RECT 51.875 0 52.375 10 ;
      RECT 51.125 0.125 51.625 9.875 ;
      RECT 50.375 0 50.875 10 ;
      RECT 49.625 0.125 50.125 9.875 ;
      RECT 48.875 0 49.375 10 ;
      RECT 48.125 0.125 48.625 9.875 ;
      RECT 47.375 0 47.875 10 ;
      RECT 46.625 0.125 47.125 9.875 ;
      RECT 45.875 0 46.375 10 ;
      RECT 45.125 0.125 45.625 9.875 ;
      RECT 44.375 0 44.875 10 ;
      RECT 43.625 0.125 44.125 9.875 ;
      RECT 42.875 0 43.375 10 ;
      RECT 42.125 0.125 42.625 9.875 ;
      RECT 41.375 0 41.875 10 ;
      RECT 40.625 0.125 41.125 9.875 ;
      RECT 39.875 0 40.375 10 ;
      RECT 39.125 0.125 39.625 9.875 ;
      RECT 38.375 0 38.875 10 ;
      RECT 37.625 0.125 38.125 9.875 ;
      RECT 36.875 0 37.375 10 ;
      RECT 36.125 0.125 36.625 9.875 ;
      RECT 35.375 0 35.875 10 ;
      RECT 34.625 0.125 35.125 9.875 ;
      RECT 33.875 0 34.375 10 ;
      RECT 33.125 0.125 33.625 9.875 ;
      RECT 32.375 0 32.875 10 ;
      RECT 31.625 0.125 32.125 9.875 ;
      RECT 30.875 0 31.375 10 ;
      RECT 30.125 0.125 30.625 9.875 ;
      RECT 29.375 0 29.875 10 ;
      RECT 28.625 0.125 29.125 9.875 ;
      RECT 27.875 0 28.375 10 ;
      RECT 27.125 0.125 27.625 9.875 ;
      RECT 26.375 0 26.875 10 ;
      RECT 25.625 0.125 26.125 9.875 ;
      RECT 24.875 0 25.375 10 ;
      RECT 24.125 0.125 24.625 9.875 ;
      RECT 23.375 0 23.875 10 ;
      RECT 22.625 0.125 23.125 9.875 ;
      RECT 21.875 0 22.375 10 ;
      RECT 21.125 0.125 21.625 9.875 ;
      RECT 20.375 0 20.875 10 ;
      RECT 19.625 0.125 20.125 9.875 ;
      RECT 18.875 0 19.375 10 ;
      RECT 18.125 0.125 18.625 9.875 ;
      RECT 17.375 0 17.875 10 ;
      RECT 16.625 0.125 17.125 9.875 ;
      RECT 15.875 0 16.375 10 ;
      RECT 15.125 0.125 15.625 9.875 ;
      RECT 14.375 0 14.875 10 ;
      RECT 13.625 0.125 14.125 9.875 ;
      RECT 12.875 0 13.375 10 ;
      RECT 12.125 0.125 12.625 9.875 ;
      RECT 11.375 0 11.875 10 ;
      RECT 10.625 0.125 11.125 9.875 ;
      RECT 9.875 0 10.375 10 ;
      RECT 9.125 0.125 9.625 9.875 ;
      RECT 8.375 0 8.875 10 ;
      RECT 7.625 0.125 8.125 9.875 ;
      RECT 6.875 0 7.375 10 ;
      RECT 6.125 0.125 6.625 9.875 ;
      RECT 5.375 0 5.875 10 ;
      RECT 4.625 0.125 5.125 9.875 ;
      RECT 3.875 0 4.375 10 ;
      RECT 3.125 0.125 3.625 9.875 ;
      RECT 2.375 0 2.875 10 ;
      RECT 1.625 0.125 2.125 9.875 ;
      RECT 0.875 0 1.375 10 ;
      RECT 0.125 0 0.625 10 ;
  END
END RIIO_EG1D80V_ESD_B2B_059x010

MACRO RIIO_HVT0D80V_CLAMP_010x230
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_HVT0D80V_CLAMP_010x230 0 0 ;
  SIZE 10 BY 230 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER C1 ;
        RECT 0.245 0.115 0.395 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 0.725 0.115 0.875 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 1.205 0.115 1.355 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 1.685 0.115 1.835 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.165 0.115 2.315 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.645 0.115 2.795 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.125 0.115 3.275 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.605 0.115 3.755 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 4.085 0.115 4.235 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.525 0.115 5.675 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.005 0.115 6.155 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.485 0.115 6.635 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.965 0.115 7.115 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.445 0.115 7.595 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.925 0.115 8.075 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.405 0.115 8.555 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.885 0.115 9.035 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.365 0.115 9.515 229.885 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER C1 ;
        RECT 0.485 0.115 0.635 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 0.965 0.115 1.115 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 1.445 0.115 1.595 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 1.925 0.115 2.075 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.405 0.115 2.555 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.885 0.115 3.035 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.365 0.115 3.515 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.845 0.115 3.995 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 4.325 0.115 4.475 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 4.805 0.115 4.955 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.285 0.115 5.435 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.765 0.115 5.915 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.245 0.115 6.395 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.725 0.115 6.875 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.205 0.115 7.355 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.685 0.115 7.835 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.165 0.115 8.315 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.645 0.115 8.795 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.125 0.115 9.275 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.605 0.115 9.755 229.885 ;
    END
  END VDD
  PIN SUB
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "sub SUB!" ;
  END SUB
  OBS
    LAYER CA ;
      RECT 0 0 10 230 ;
    LAYER M1 ;
      RECT 0 0 10 230 ;
    LAYER V1 ;
      RECT 0 0 10 230 ;
    LAYER M2 ;
      RECT 0 0 10 230 ;
    LAYER CB ;
      RECT 0 0 10 230 ;
    LAYER AY ;
      RECT 0 0 10 230 ;
    LAYER C1 ;
      RECT 9.605 0.115 9.755 229.885 ;
      RECT 9.365 0.115 9.515 229.885 ;
      RECT 9.125 0.115 9.275 229.885 ;
      RECT 8.885 0.115 9.035 229.885 ;
      RECT 8.645 0.115 8.795 229.885 ;
      RECT 8.405 0.115 8.555 229.885 ;
      RECT 8.165 0.115 8.315 229.885 ;
      RECT 7.925 0.115 8.075 229.885 ;
      RECT 7.685 0.115 7.835 229.885 ;
      RECT 7.445 0.115 7.595 229.885 ;
      RECT 7.205 0.115 7.355 229.885 ;
      RECT 6.965 0.115 7.115 229.885 ;
      RECT 6.725 0.115 6.875 229.885 ;
      RECT 6.485 0.115 6.635 229.885 ;
      RECT 6.245 0.115 6.395 229.885 ;
      RECT 6.005 0.115 6.155 229.885 ;
      RECT 5.765 0.115 5.915 229.885 ;
      RECT 5.525 0.115 5.675 229.885 ;
      RECT 5.285 0.115 5.435 229.885 ;
      RECT 5.045 0.628 5.195 182.428 ;
      RECT 5.045 182.731 5.195 229.885 ;
      RECT 4.805 0.115 4.955 229.885 ;
      RECT 4.565 0.628 4.715 182.428 ;
      RECT 4.565 182.731 4.715 229.885 ;
      RECT 4.325 0.115 4.475 229.885 ;
      RECT 4.085 0.115 4.235 229.885 ;
      RECT 3.845 0.115 3.995 229.885 ;
      RECT 3.605 0.115 3.755 229.885 ;
      RECT 3.365 0.115 3.515 229.885 ;
      RECT 3.125 0.115 3.275 229.885 ;
      RECT 2.885 0.115 3.035 229.885 ;
      RECT 2.645 0.115 2.795 229.885 ;
      RECT 2.405 0.115 2.555 229.885 ;
      RECT 2.165 0.115 2.315 229.885 ;
      RECT 1.925 0.115 2.075 229.885 ;
      RECT 1.685 0.115 1.835 229.885 ;
      RECT 1.445 0.115 1.595 229.885 ;
      RECT 1.205 0.115 1.355 229.885 ;
      RECT 0.965 0.115 1.115 229.885 ;
      RECT 0.725 0.115 0.875 229.885 ;
      RECT 0.485 0.115 0.635 229.885 ;
      RECT 0.245 0.115 0.395 229.885 ;
  END
END RIIO_HVT0D80V_CLAMP_010x230

MACRO RIIO_HVT0D80V_CLAMP_059x057
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_HVT0D80V_CLAMP_059x057 0 0 ;
  SIZE 59.25 BY 57.28 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER C1 ;
        RECT 0.875 0 1.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.375 0 2.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.875 0 4.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.375 0 5.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.875 0 7.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.375 0 8.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.875 0 10.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 11.375 0 11.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 12.875 0 13.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 14.375 0 14.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 15.875 0 16.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 17.375 0 17.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 18.875 0 19.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 20.375 0 20.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 21.875 0 22.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 23.375 0 23.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 24.875 0 25.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 26.375 0 26.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 27.875 0 28.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 29.375 0 29.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 30.875 0 31.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 32.375 0 32.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 33.875 0 34.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 35.375 0 35.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 36.875 0 37.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 38.375 0 38.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 39.875 0 40.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 41.375 0 41.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 42.875 0 43.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 44.375 0 44.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 45.875 0 46.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 47.375 0 47.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 48.875 0 49.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 50.375 0 50.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 51.875 0 52.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 53.375 0 53.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 54.875 0 55.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 56.375 0 56.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 57.875 0 58.375 57.28 ;
    END
  END VSS
  PIN SUB
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "sub SUB!" ;
    PORT
      LAYER C1 ;
        RECT 0.125 0 0.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 58.625 0 59.125 57.28 ;
    END
  END SUB
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER C1 ;
        RECT 1.625 0 2.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.125 0 3.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 4.625 0 5.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.125 0 6.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.625 0 8.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.125 0 9.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 10.625 0 11.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 12.125 0 12.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 13.625 0 14.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 15.125 0 15.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 16.625 0 17.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 18.125 0 18.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 19.625 0 20.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 21.125 0 21.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 22.625 0 23.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 24.125 0 24.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 25.625 0 26.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 27.125 0 27.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 28.625 0 29.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 30.125 0 30.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 31.625 0 32.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 33.125 0 33.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 34.625 0 35.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 36.125 0 36.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 37.625 0 38.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 39.125 0 39.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 40.625 0 41.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 42.125 0 42.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 43.625 0 44.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 45.125 0 45.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 46.625 0 47.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 48.125 0 48.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 49.625 0 50.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 51.125 0 51.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 52.625 0 53.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 54.125 0 54.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 55.625 0 56.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 57.125 0 57.625 57.28 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 59.25 57.28 ;
    LAYER M1 ;
      RECT 0 0 59.25 57.28 ;
    LAYER V1 ;
      RECT 0 0 59.25 57.28 ;
    LAYER M2 ;
      RECT 0 0 59.25 57.28 ;
    LAYER CB ;
      RECT 0 0 59.25 57.28 ;
    LAYER AY ;
      RECT 0 0 59.25 57.28 ;
    LAYER C1 ;
      RECT 58.625 0 59.125 57.28 ;
      RECT 57.875 0 58.375 57.28 ;
      RECT 57.125 0 57.625 57.28 ;
      RECT 56.375 0 56.875 57.28 ;
      RECT 55.625 0 56.125 57.28 ;
      RECT 54.875 0 55.375 57.28 ;
      RECT 54.125 0 54.625 57.28 ;
      RECT 53.375 0 53.875 57.28 ;
      RECT 52.625 0 53.125 57.28 ;
      RECT 51.875 0 52.375 57.28 ;
      RECT 51.125 0 51.625 57.28 ;
      RECT 50.375 0 50.875 57.28 ;
      RECT 49.625 0 50.125 57.28 ;
      RECT 48.875 0 49.375 57.28 ;
      RECT 48.125 0 48.625 57.28 ;
      RECT 47.375 0 47.875 57.28 ;
      RECT 46.625 0 47.125 57.28 ;
      RECT 45.875 0 46.375 57.28 ;
      RECT 45.125 0 45.625 57.28 ;
      RECT 44.375 0 44.875 57.28 ;
      RECT 43.625 0 44.125 57.28 ;
      RECT 42.875 0 43.375 57.28 ;
      RECT 42.125 0 42.625 57.28 ;
      RECT 41.375 0 41.875 57.28 ;
      RECT 40.625 0 41.125 57.28 ;
      RECT 39.875 0 40.375 57.28 ;
      RECT 39.125 0 39.625 57.28 ;
      RECT 38.375 0 38.875 57.28 ;
      RECT 37.625 0 38.125 57.28 ;
      RECT 36.875 0 37.375 57.28 ;
      RECT 36.125 0 36.625 57.28 ;
      RECT 35.375 0 35.875 57.28 ;
      RECT 34.625 0 35.125 57.28 ;
      RECT 33.875 0 34.375 57.28 ;
      RECT 33.125 0 33.625 57.28 ;
      RECT 32.375 0 32.875 57.28 ;
      RECT 31.625 0 32.125 57.28 ;
      RECT 30.875 0 31.375 57.28 ;
      RECT 30.125 0 30.625 57.28 ;
      RECT 29.375 0 29.875 57.28 ;
      RECT 28.625 0 29.125 57.28 ;
      RECT 27.875 0 28.375 57.28 ;
      RECT 27.125 0 27.625 57.28 ;
      RECT 26.375 0 26.875 57.28 ;
      RECT 25.625 0 26.125 57.28 ;
      RECT 24.875 0 25.375 57.28 ;
      RECT 24.125 0 24.625 57.28 ;
      RECT 23.375 0 23.875 57.28 ;
      RECT 22.625 0 23.125 57.28 ;
      RECT 21.875 0 22.375 57.28 ;
      RECT 21.125 0 21.625 57.28 ;
      RECT 20.375 0 20.875 57.28 ;
      RECT 19.625 0 20.125 57.28 ;
      RECT 18.875 0 19.375 57.28 ;
      RECT 18.125 0 18.625 57.28 ;
      RECT 17.375 0 17.875 57.28 ;
      RECT 16.625 0 17.125 57.28 ;
      RECT 15.875 0 16.375 57.28 ;
      RECT 15.125 0 15.625 57.28 ;
      RECT 14.375 0 14.875 57.28 ;
      RECT 13.625 0 14.125 57.28 ;
      RECT 12.875 0 13.375 57.28 ;
      RECT 12.125 0 12.625 57.28 ;
      RECT 11.375 0 11.875 57.28 ;
      RECT 10.625 0 11.125 57.28 ;
      RECT 9.875 0 10.375 57.28 ;
      RECT 9.125 0 9.625 57.28 ;
      RECT 8.375 0 8.875 57.28 ;
      RECT 7.625 0 8.125 57.28 ;
      RECT 6.875 0 7.375 57.28 ;
      RECT 6.125 0 6.625 57.28 ;
      RECT 5.375 0 5.875 57.28 ;
      RECT 4.625 0 5.125 57.28 ;
      RECT 3.875 0 4.375 57.28 ;
      RECT 3.125 0 3.625 57.28 ;
      RECT 2.375 0 2.875 57.28 ;
      RECT 1.625 0 2.125 57.28 ;
      RECT 0.875 0 1.375 57.28 ;
      RECT 0.125 0 0.625 57.28 ;
  END
END RIIO_HVT0D80V_CLAMP_059x057

MACRO RIIO_RVT0D80V_CLAMP_010x230
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_RVT0D80V_CLAMP_010x230 0 0 ;
  SIZE 10 BY 230 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER C1 ;
        RECT 0.245 0.115 0.395 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 0.725 0.115 0.875 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 1.205 0.115 1.355 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 1.685 0.115 1.835 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.165 0.115 2.315 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.645 0.115 2.795 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.125 0.115 3.275 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.605 0.115 3.755 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 4.085 0.115 4.235 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.525 0.115 5.675 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.005 0.115 6.155 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.485 0.115 6.635 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.965 0.115 7.115 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.445 0.115 7.595 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.925 0.115 8.075 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.405 0.115 8.555 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.885 0.115 9.035 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.365 0.115 9.515 229.885 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER C1 ;
        RECT 0.485 0.115 0.635 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 0.965 0.115 1.115 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 1.445 0.115 1.595 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 1.925 0.115 2.075 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.405 0.115 2.555 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.885 0.115 3.035 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.365 0.115 3.515 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.845 0.115 3.995 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 4.325 0.115 4.475 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 4.805 0.115 4.955 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.285 0.115 5.435 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.765 0.115 5.915 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.245 0.115 6.395 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.725 0.115 6.875 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.205 0.115 7.355 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.685 0.115 7.835 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.165 0.115 8.315 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.645 0.115 8.795 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.125 0.115 9.275 229.885 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.605 0.115 9.755 229.885 ;
    END
  END VDD
  PIN SUB
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "sub SUB!" ;
  END SUB
  OBS
    LAYER CA ;
      RECT 0 0 10 230 ;
    LAYER M1 ;
      RECT 0 0 10 230 ;
    LAYER V1 ;
      RECT 0 0 10 230 ;
    LAYER M2 ;
      RECT 0 0 10 230 ;
    LAYER CB ;
      RECT 0 0 10 230 ;
    LAYER AY ;
      RECT 0 0 10 230 ;
    LAYER C1 ;
      RECT 9.605 0.115 9.755 229.885 ;
      RECT 9.365 0.115 9.515 229.885 ;
      RECT 9.125 0.115 9.275 229.885 ;
      RECT 8.885 0.115 9.035 229.885 ;
      RECT 8.645 0.115 8.795 229.885 ;
      RECT 8.405 0.115 8.555 229.885 ;
      RECT 8.165 0.115 8.315 229.885 ;
      RECT 7.925 0.115 8.075 229.885 ;
      RECT 7.685 0.115 7.835 229.885 ;
      RECT 7.445 0.115 7.595 229.885 ;
      RECT 7.205 0.115 7.355 229.885 ;
      RECT 6.965 0.115 7.115 229.885 ;
      RECT 6.725 0.115 6.875 229.885 ;
      RECT 6.485 0.115 6.635 229.885 ;
      RECT 6.245 0.115 6.395 229.885 ;
      RECT 6.005 0.115 6.155 229.885 ;
      RECT 5.765 0.115 5.915 229.885 ;
      RECT 5.525 0.115 5.675 229.885 ;
      RECT 5.285 0.115 5.435 229.885 ;
      RECT 5.045 0.628 5.195 182.428 ;
      RECT 5.045 182.731 5.195 229.885 ;
      RECT 4.805 0.115 4.955 229.885 ;
      RECT 4.565 0.628 4.715 182.428 ;
      RECT 4.565 182.731 4.715 229.885 ;
      RECT 4.325 0.115 4.475 229.885 ;
      RECT 4.085 0.115 4.235 229.885 ;
      RECT 3.845 0.115 3.995 229.885 ;
      RECT 3.605 0.115 3.755 229.885 ;
      RECT 3.365 0.115 3.515 229.885 ;
      RECT 3.125 0.115 3.275 229.885 ;
      RECT 2.885 0.115 3.035 229.885 ;
      RECT 2.645 0.115 2.795 229.885 ;
      RECT 2.405 0.115 2.555 229.885 ;
      RECT 2.165 0.115 2.315 229.885 ;
      RECT 1.925 0.115 2.075 229.885 ;
      RECT 1.685 0.115 1.835 229.885 ;
      RECT 1.445 0.115 1.595 229.885 ;
      RECT 1.205 0.115 1.355 229.885 ;
      RECT 0.965 0.115 1.115 229.885 ;
      RECT 0.725 0.115 0.875 229.885 ;
      RECT 0.485 0.115 0.635 229.885 ;
      RECT 0.245 0.115 0.395 229.885 ;
  END
END RIIO_RVT0D80V_CLAMP_010x230

MACRO RIIO_RVT0D80V_CLAMP_059x057
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_RVT0D80V_CLAMP_059x057 0 0 ;
  SIZE 59.25 BY 57.28 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER C1 ;
        RECT 0.875 0 1.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 2.375 0 2.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.875 0 4.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 5.375 0 5.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.875 0 7.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 8.375 0 8.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.875 0 10.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 11.375 0 11.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 12.875 0 13.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 14.375 0 14.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 15.875 0 16.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 17.375 0 17.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 18.875 0 19.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 20.375 0 20.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 21.875 0 22.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 23.375 0 23.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 24.875 0 25.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 26.375 0 26.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 27.875 0 28.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 29.375 0 29.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 30.875 0 31.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 32.375 0 32.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 33.875 0 34.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 35.375 0 35.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 36.875 0 37.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 38.375 0 38.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 39.875 0 40.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 41.375 0 41.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 42.875 0 43.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 44.375 0 44.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 45.875 0 46.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 47.375 0 47.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 48.875 0 49.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 50.375 0 50.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 51.875 0 52.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 53.375 0 53.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 54.875 0 55.375 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 56.375 0 56.875 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 57.875 0 58.375 57.28 ;
    END
  END VSS
  PIN SUB
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "sub SUB!" ;
    PORT
      LAYER C1 ;
        RECT 0.125 0 0.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 58.625 0 59.125 57.28 ;
    END
  END SUB
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER C1 ;
        RECT 1.625 0 2.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 3.125 0 3.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 4.625 0 5.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 6.125 0 6.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 7.625 0 8.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 9.125 0 9.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 10.625 0 11.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 12.125 0 12.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 13.625 0 14.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 15.125 0 15.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 16.625 0 17.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 18.125 0 18.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 19.625 0 20.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 21.125 0 21.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 22.625 0 23.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 24.125 0 24.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 25.625 0 26.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 27.125 0 27.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 28.625 0 29.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 30.125 0 30.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 31.625 0 32.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 33.125 0 33.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 34.625 0 35.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 36.125 0 36.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 37.625 0 38.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 39.125 0 39.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 40.625 0 41.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 42.125 0 42.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 43.625 0 44.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 45.125 0 45.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 46.625 0 47.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 48.125 0 48.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 49.625 0 50.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 51.125 0 51.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 52.625 0 53.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 54.125 0 54.625 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 55.625 0 56.125 57.28 ;
    END
    PORT
      LAYER C1 ;
        RECT 57.125 0 57.625 57.28 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 59.25 57.28 ;
    LAYER M1 ;
      RECT 0 0 59.25 57.28 ;
    LAYER V1 ;
      RECT 0 0 59.25 57.28 ;
    LAYER M2 ;
      RECT 0 0 59.25 57.28 ;
    LAYER CB ;
      RECT 0 0 59.25 57.28 ;
    LAYER AY ;
      RECT 0 0 59.25 57.28 ;
    LAYER C1 ;
      RECT 58.625 0 59.125 57.28 ;
      RECT 57.875 0 58.375 57.28 ;
      RECT 57.125 0 57.625 57.28 ;
      RECT 56.375 0 56.875 57.28 ;
      RECT 55.625 0 56.125 57.28 ;
      RECT 54.875 0 55.375 57.28 ;
      RECT 54.125 0 54.625 57.28 ;
      RECT 53.375 0 53.875 57.28 ;
      RECT 52.625 0 53.125 57.28 ;
      RECT 51.875 0 52.375 57.28 ;
      RECT 51.125 0 51.625 57.28 ;
      RECT 50.375 0 50.875 57.28 ;
      RECT 49.625 0 50.125 57.28 ;
      RECT 48.875 0 49.375 57.28 ;
      RECT 48.125 0 48.625 57.28 ;
      RECT 47.375 0 47.875 57.28 ;
      RECT 46.625 0 47.125 57.28 ;
      RECT 45.875 0 46.375 57.28 ;
      RECT 45.125 0 45.625 57.28 ;
      RECT 44.375 0 44.875 57.28 ;
      RECT 43.625 0 44.125 57.28 ;
      RECT 42.875 0 43.375 57.28 ;
      RECT 42.125 0 42.625 57.28 ;
      RECT 41.375 0 41.875 57.28 ;
      RECT 40.625 0 41.125 57.28 ;
      RECT 39.875 0 40.375 57.28 ;
      RECT 39.125 0 39.625 57.28 ;
      RECT 38.375 0 38.875 57.28 ;
      RECT 37.625 0 38.125 57.28 ;
      RECT 36.875 0 37.375 57.28 ;
      RECT 36.125 0 36.625 57.28 ;
      RECT 35.375 0 35.875 57.28 ;
      RECT 34.625 0 35.125 57.28 ;
      RECT 33.875 0 34.375 57.28 ;
      RECT 33.125 0 33.625 57.28 ;
      RECT 32.375 0 32.875 57.28 ;
      RECT 31.625 0 32.125 57.28 ;
      RECT 30.875 0 31.375 57.28 ;
      RECT 30.125 0 30.625 57.28 ;
      RECT 29.375 0 29.875 57.28 ;
      RECT 28.625 0 29.125 57.28 ;
      RECT 27.875 0 28.375 57.28 ;
      RECT 27.125 0 27.625 57.28 ;
      RECT 26.375 0 26.875 57.28 ;
      RECT 25.625 0 26.125 57.28 ;
      RECT 24.875 0 25.375 57.28 ;
      RECT 24.125 0 24.625 57.28 ;
      RECT 23.375 0 23.875 57.28 ;
      RECT 22.625 0 23.125 57.28 ;
      RECT 21.875 0 22.375 57.28 ;
      RECT 21.125 0 21.625 57.28 ;
      RECT 20.375 0 20.875 57.28 ;
      RECT 19.625 0 20.125 57.28 ;
      RECT 18.875 0 19.375 57.28 ;
      RECT 18.125 0 18.625 57.28 ;
      RECT 17.375 0 17.875 57.28 ;
      RECT 16.625 0 17.125 57.28 ;
      RECT 15.875 0 16.375 57.28 ;
      RECT 15.125 0 15.625 57.28 ;
      RECT 14.375 0 14.875 57.28 ;
      RECT 13.625 0 14.125 57.28 ;
      RECT 12.875 0 13.375 57.28 ;
      RECT 12.125 0 12.625 57.28 ;
      RECT 11.375 0 11.875 57.28 ;
      RECT 10.625 0 11.125 57.28 ;
      RECT 9.875 0 10.375 57.28 ;
      RECT 9.125 0 9.625 57.28 ;
      RECT 8.375 0 8.875 57.28 ;
      RECT 7.625 0 8.125 57.28 ;
      RECT 6.875 0 7.375 57.28 ;
      RECT 6.125 0 6.625 57.28 ;
      RECT 5.375 0 5.875 57.28 ;
      RECT 4.625 0 5.125 57.28 ;
      RECT 3.875 0 4.375 57.28 ;
      RECT 3.125 0 3.625 57.28 ;
      RECT 2.375 0 2.875 57.28 ;
      RECT 1.625 0 2.125 57.28 ;
      RECT 0.875 0 1.375 57.28 ;
      RECT 0.125 0 0.625 57.28 ;
  END
END RIIO_RVT0D80V_CLAMP_059x057

MACRO RIIO_RVT36G1_RESETGEN16
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_RVT36G1_RESETGEN16 0 0 ;
  SIZE 25.172 BY 5.16 ;
  SYMMETRY X Y ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER M2 ;
        RECT 0 0 25.172 0.12 ;
      LAYER C1 ;
        RECT 24.996 0 25.136 5.16 ;
        RECT 24.476 0 24.616 5.16 ;
        RECT 21.356 0 21.496 5.16 ;
        RECT 20.836 0 20.976 2.16 ;
        RECT 20.316 0 20.456 5.16 ;
        RECT 19.276 0 19.416 5.16 ;
        RECT 18.756 0 18.896 5.16 ;
        RECT 17.716 0 17.856 5.16 ;
        RECT 17.196 0 17.336 5.16 ;
        RECT 16.676 0 16.816 5.16 ;
        RECT 16.156 0 16.296 5.16 ;
        RECT 15.636 0 15.776 5.16 ;
        RECT 14.596 0 14.736 5.16 ;
        RECT 14.076 0 14.216 5.16 ;
        RECT 13.036 0 13.176 5.16 ;
        RECT 12.516 0 12.656 5.16 ;
        RECT 11.996 0 12.136 5.16 ;
        RECT 11.476 0 11.616 5.16 ;
        RECT 10.956 0 11.096 5.16 ;
        RECT 10.436 0 10.576 5.16 ;
        RECT 9.916 0 10.056 5.16 ;
        RECT 9.396 0 9.536 5.16 ;
        RECT 7.836 0 7.976 5.16 ;
        RECT 6.796 0 6.936 5.16 ;
        RECT 5.756 0 5.896 5.16 ;
        RECT 5.236 0 5.376 5.16 ;
        RECT 3.676 0 3.816 5.16 ;
        RECT 2.116 0 2.256 5.16 ;
        RECT 1.596 0 1.736 5.16 ;
    END
  END VDD
  PIN TIMER_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.642857 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 7.316 0 7.456 5.16 ;
    END
  END TIMER_I[7]
  PIN TIMER_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.092262 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 15.116 0 15.256 5.16 ;
    END
  END TIMER_I[6]
  PIN TIMER_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.092262 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.796 0 19.936 5.16 ;
    END
  END TIMER_I[5]
  PIN TIMER_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 6.654762 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 24.216 0 24.356 5.16 ;
    END
  END TIMER_I[4]
  PIN TIMER_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8e-05 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.64881 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 18.236 0 18.376 5.16 ;
    END
  END TIMER_I[3]
  PIN TIMER_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.514881 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 13.556 0 13.696 5.16 ;
    END
  END TIMER_I[2]
  PIN TIMER_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.071429 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 8.876 0 9.016 5.16 ;
    END
  END TIMER_I[1]
  PIN TIMER_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 3.473214 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.716 0 4.856 5.16 ;
    END
  END TIMER_I[0]
  PIN RES_N_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 4.75 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 0.816 0 0.956 5.16 ;
    END
  END RES_N_I[3]
  PIN RES_N_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 5.077381 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 0.556 0 0.696 5.16 ;
    END
  END RES_N_I[2]
  PIN RES_N_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 6.72619 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 0.296 0 0.436 5.16 ;
    END
  END RES_N_I[1]
  PIN RES_N_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 6.696429 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 0.036 0 0.176 5.16 ;
    END
  END RES_N_I[0]
  PIN RESET_N_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16896 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.196 0 4.336 5.16 ;
    END
  END RESET_N_O
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER M2 ;
        RECT 0 0.24 25.172 0.36 ;
      LAYER C1 ;
        RECT 24.736 0 24.876 5.16 ;
        RECT 23.176 0 23.316 5.16 ;
        RECT 22.656 0 22.796 5.16 ;
        RECT 22.136 0 22.276 5.16 ;
        RECT 21.616 0 21.756 5.16 ;
        RECT 21.096 0 21.236 5.16 ;
        RECT 20.576 0 20.716 5.16 ;
        RECT 20.056 0 20.196 5.16 ;
        RECT 19.536 0 19.676 5.16 ;
        RECT 19.016 0 19.156 5.16 ;
        RECT 18.496 0 18.636 5.16 ;
        RECT 17.976 0 18.116 5.16 ;
        RECT 17.456 0 17.596 5.16 ;
        RECT 16.936 0 17.076 5.16 ;
        RECT 16.416 0 16.556 5.16 ;
        RECT 15.896 0 16.036 5.16 ;
        RECT 15.376 0 15.516 5.16 ;
        RECT 14.856 0 14.996 5.16 ;
        RECT 14.336 0 14.476 5.16 ;
        RECT 13.816 0 13.956 5.16 ;
        RECT 13.296 0 13.436 5.16 ;
        RECT 12.776 0 12.916 5.16 ;
        RECT 12.256 0 12.396 5.16 ;
        RECT 11.736 0 11.876 5.16 ;
        RECT 11.216 0 11.356 5.16 ;
        RECT 10.696 0 10.836 5.16 ;
        RECT 10.176 0 10.316 5.16 ;
        RECT 9.656 0 9.796 5.16 ;
        RECT 9.136 0 9.276 5.16 ;
        RECT 8.616 0 8.756 5.16 ;
        RECT 8.096 0 8.236 5.16 ;
        RECT 7.576 0 7.716 5.16 ;
        RECT 7.056 0 7.196 5.16 ;
        RECT 6.536 0 6.676 5.16 ;
        RECT 6.016 0 6.156 5.16 ;
        RECT 5.496 0 5.636 5.16 ;
        RECT 4.976 0 5.116 5.16 ;
        RECT 4.456 0 4.596 5.16 ;
        RECT 3.936 0 4.076 5.16 ;
        RECT 3.416 0 3.556 5.16 ;
        RECT 2.896 0 3.036 5.16 ;
        RECT 2.376 0 2.516 5.16 ;
        RECT 1.856 0 1.996 5.16 ;
        RECT 1.336 0 1.476 5.16 ;
    END
  END VSS
  PIN EN_N_CS_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 9.464286 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.956 0 24.096 5.16 ;
    END
  END EN_N_CS_I
  PIN CLK_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16192 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 22.916 0 23.056 5.16 ;
    END
  END CLK_O
  PIN EN_N_CR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 6.446429 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.696 0 23.836 5.16 ;
    END
  END EN_N_CR_I
  OBS
    LAYER CA ;
      RECT 0 0 25.172 5.16 ;
    LAYER M1 ;
      RECT 0 0 25.172 5.16 ;
    LAYER V1 ;
      RECT 0 0 25.172 5.16 ;
    LAYER M2 ;
      RECT 0 0 25.172 5.16 ;
    LAYER CB ;
      RECT 0 0 25.172 5.16 ;
    LAYER AY ;
      RECT 0 0 25.172 5.16 ;
    LAYER C1 ;
      RECT 18.236 0 18.376 5.16 ;
      RECT 18.235 1.82 18.376 1.9 ;
      RECT 24.996 0 25.136 5.16 ;
      RECT 24.736 0 24.876 5.16 ;
      RECT 24.476 0 24.616 5.16 ;
      RECT 24.216 0 24.356 5.16 ;
      RECT 23.956 0 24.096 5.16 ;
      RECT 23.696 0 23.836 5.16 ;
      RECT 23.436 0 23.576 0.72 ;
      RECT 23.436 0.84 23.576 3.6 ;
      RECT 23.436 3.72 23.576 5.16 ;
      RECT 23.176 0 23.316 5.16 ;
      RECT 22.916 0 23.056 5.16 ;
      RECT 22.656 0 22.796 5.16 ;
      RECT 22.396 0 22.536 0.72 ;
      RECT 22.396 0.84 22.536 2.16 ;
      RECT 22.396 2.28 22.536 3.6 ;
      RECT 22.396 3.72 22.536 5.16 ;
      RECT 22.136 0 22.276 5.16 ;
      RECT 21.876 0 22.016 0.72 ;
      RECT 21.876 0.84 22.016 2.16 ;
      RECT 21.876 2.28 22.016 4.32 ;
      RECT 21.876 4.44 22.016 5.16 ;
      RECT 21.616 0 21.756 5.16 ;
      RECT 21.356 0 21.496 5.16 ;
      RECT 21.096 0 21.236 5.16 ;
      RECT 20.836 0 20.976 2.16 ;
      RECT 20.836 2.28 20.976 2.62 ;
      RECT 20.836 2.7 20.976 3.6 ;
      RECT 20.836 3.72 20.976 5.16 ;
      RECT 20.576 0 20.716 5.16 ;
      RECT 20.316 0 20.456 5.16 ;
      RECT 20.056 0 20.196 5.16 ;
      RECT 19.796 0 19.936 5.16 ;
      RECT 19.536 0 19.676 5.16 ;
      RECT 19.276 0 19.416 5.16 ;
      RECT 19.016 0 19.156 5.16 ;
      RECT 18.756 0 18.896 5.16 ;
      RECT 18.496 0 18.636 5.16 ;
      RECT 17.976 0 18.116 5.16 ;
      RECT 17.716 0 17.856 5.16 ;
      RECT 17.456 0 17.596 5.16 ;
      RECT 17.196 0 17.336 5.16 ;
      RECT 16.936 0 17.076 5.16 ;
      RECT 16.676 0 16.816 5.16 ;
      RECT 16.416 0 16.556 5.16 ;
      RECT 16.156 0 16.296 5.16 ;
      RECT 15.896 0 16.036 5.16 ;
      RECT 15.636 0 15.776 5.16 ;
      RECT 15.376 0 15.516 5.16 ;
      RECT 15.116 0 15.256 5.16 ;
      RECT 14.856 0 14.996 5.16 ;
      RECT 14.596 0 14.736 5.16 ;
      RECT 14.336 0 14.476 5.16 ;
      RECT 14.076 0 14.216 5.16 ;
      RECT 13.816 0 13.956 5.16 ;
      RECT 13.556 0 13.696 5.16 ;
      RECT 13.296 0 13.436 5.16 ;
      RECT 13.036 0 13.176 5.16 ;
      RECT 12.776 0 12.916 5.16 ;
      RECT 12.516 0 12.656 5.16 ;
      RECT 12.256 0 12.396 5.16 ;
      RECT 11.996 0 12.136 5.16 ;
      RECT 11.736 0 11.876 5.16 ;
      RECT 11.476 0 11.616 5.16 ;
      RECT 11.216 0 11.356 5.16 ;
      RECT 10.956 0 11.096 5.16 ;
      RECT 10.696 0 10.836 5.16 ;
      RECT 10.436 0 10.576 5.16 ;
      RECT 10.176 0 10.316 5.16 ;
      RECT 9.916 0 10.056 5.16 ;
      RECT 9.656 0 9.796 5.16 ;
      RECT 9.396 0 9.536 5.16 ;
      RECT 9.136 0 9.276 5.16 ;
      RECT 8.876 0 9.016 5.16 ;
      RECT 8.616 0 8.756 5.16 ;
      RECT 8.356 0 8.496 0.72 ;
      RECT 8.356 0.84 8.496 1.44 ;
      RECT 8.356 1.56 8.496 5.16 ;
      RECT 8.096 0 8.236 5.16 ;
      RECT 7.836 0 7.976 5.16 ;
      RECT 7.576 0 7.716 5.16 ;
      RECT 7.316 0 7.456 5.16 ;
      RECT 7.056 0 7.196 5.16 ;
      RECT 6.796 0 6.936 5.16 ;
      RECT 6.536 0 6.676 5.16 ;
      RECT 6.276 0 6.416 0.72 ;
      RECT 6.276 0.84 6.416 3.6 ;
      RECT 6.276 3.72 6.416 5.16 ;
      RECT 6.016 0 6.156 5.16 ;
      RECT 5.756 0 5.896 5.16 ;
      RECT 5.496 0 5.636 5.16 ;
      RECT 5.236 0 5.376 5.16 ;
      RECT 4.976 0 5.116 5.16 ;
      RECT 4.716 0 4.856 5.16 ;
      RECT 4.456 0 4.596 5.16 ;
      RECT 4.196 0 4.336 5.16 ;
      RECT 3.936 0 4.076 5.16 ;
      RECT 3.676 0 3.816 5.16 ;
      RECT 3.416 0 3.556 5.16 ;
      RECT 3.156 0 3.296 1.44 ;
      RECT 3.156 1.56 3.296 2.88 ;
      RECT 3.156 3 3.296 5.16 ;
      RECT 2.896 0 3.036 5.16 ;
      RECT 2.636 0 2.776 0.72 ;
      RECT 2.636 0.84 2.776 2.88 ;
      RECT 2.636 3 2.776 4.32 ;
      RECT 2.636 4.44 2.776 5.16 ;
      RECT 2.376 0 2.516 5.16 ;
      RECT 2.116 0 2.256 5.16 ;
      RECT 1.856 0 1.996 5.16 ;
      RECT 1.596 0 1.736 5.16 ;
      RECT 1.336 0 1.476 5.16 ;
      RECT 1.076 0 1.216 1.44 ;
      RECT 1.076 1.56 1.216 2.88 ;
      RECT 1.076 3 1.216 5.16 ;
      RECT 0.816 0 0.956 5.16 ;
      RECT 0.556 0 0.696 5.16 ;
      RECT 0.296 0 0.436 5.16 ;
      RECT 0.036 0 0.176 5.16 ;
  END
END RIIO_RVT36G1_RESETGEN16

MACRO RIIO_RVT36G1_RESETGEN27
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_RVT36G1_RESETGEN27 0 0 ;
  SIZE 25.172 BY 6.6 ;
  SYMMETRY X Y ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER M2 ;
        RECT 0 0 25.172 0.12 ;
      LAYER C1 ;
        RECT 24.996 0 25.136 6.6 ;
        RECT 24.476 0 24.616 6.6 ;
        RECT 21.356 0 21.496 6.6 ;
        RECT 20.836 0 20.976 2.16 ;
        RECT 20.316 0 20.456 6.6 ;
        RECT 19.276 0 19.416 6.6 ;
        RECT 18.756 0 18.896 6.6 ;
        RECT 17.716 0 17.856 6.6 ;
        RECT 17.196 0 17.336 6.6 ;
        RECT 16.676 0 16.816 6.6 ;
        RECT 16.156 0 16.296 6.6 ;
        RECT 15.636 0 15.776 6.6 ;
        RECT 14.596 0 14.736 6.6 ;
        RECT 14.076 0 14.216 6.6 ;
        RECT 13.036 0 13.176 6.6 ;
        RECT 12.516 0 12.656 6.6 ;
        RECT 11.996 0 12.136 6.6 ;
        RECT 11.476 0 11.616 6.6 ;
        RECT 10.956 0 11.096 6.6 ;
        RECT 10.436 0 10.576 6.6 ;
        RECT 9.916 0 10.056 6.6 ;
        RECT 9.396 0 9.536 6.6 ;
        RECT 7.836 0 7.976 6.6 ;
        RECT 6.796 0 6.936 6.6 ;
        RECT 5.756 0 5.896 6.6 ;
        RECT 5.236 0 5.376 6.6 ;
        RECT 3.676 0 3.816 6.6 ;
        RECT 2.116 0 2.256 6.6 ;
        RECT 1.596 0 1.736 6.6 ;
    END
  END VDD
  PIN TIMER_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.642857 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 7.316 0 7.456 6.6 ;
    END
  END TIMER_I[7]
  PIN TIMER_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.092262 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 15.116 0 15.256 6.6 ;
    END
  END TIMER_I[6]
  PIN TIMER_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.092262 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.796 0 19.936 6.6 ;
    END
  END TIMER_I[5]
  PIN TIMER_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 6.654762 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 24.216 0 24.356 6.6 ;
    END
  END TIMER_I[4]
  PIN TIMER_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8e-05 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.64881 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 18.236 0 18.376 6.6 ;
    END
  END TIMER_I[3]
  PIN TIMER_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.514881 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 13.556 0 13.696 6.6 ;
    END
  END TIMER_I[2]
  PIN TIMER_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 2.071429 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 8.876 0 9.016 6.6 ;
    END
  END TIMER_I[1]
  PIN TIMER_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 3.473214 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.716 0 4.856 6.6 ;
    END
  END TIMER_I[0]
  PIN RES_N_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 4.75 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 0.816 0 0.956 6.6 ;
    END
  END RES_N_I[3]
  PIN RES_N_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 5.077381 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 0.556 0 0.696 6.6 ;
    END
  END RES_N_I[2]
  PIN RES_N_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 6.72619 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 0.296 0 0.436 6.6 ;
    END
  END RES_N_I[1]
  PIN RES_N_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01344 LAYER C1 ;
      ANTENNAMAXAREACAR 6.696429 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 0.036 0 0.176 6.6 ;
    END
  END RES_N_I[0]
  PIN RESET_N_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16896 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.196 0 4.336 6.6 ;
    END
  END RESET_N_O
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER M2 ;
        RECT 0 0.24 25.172 0.36 ;
      LAYER C1 ;
        RECT 24.736 0 24.876 6.6 ;
        RECT 23.176 0 23.316 6.6 ;
        RECT 22.656 0 22.796 6.6 ;
        RECT 22.136 0 22.276 6.6 ;
        RECT 21.616 0 21.756 6.6 ;
        RECT 21.096 0 21.236 6.6 ;
        RECT 20.576 0 20.716 6.6 ;
        RECT 20.056 0 20.196 6.6 ;
        RECT 19.536 0 19.676 6.6 ;
        RECT 19.016 0 19.156 6.6 ;
        RECT 18.496 0 18.636 6.6 ;
        RECT 17.976 0 18.116 6.6 ;
        RECT 17.456 0 17.596 6.6 ;
        RECT 16.936 0 17.076 6.6 ;
        RECT 16.416 0 16.556 6.6 ;
        RECT 15.896 0 16.036 6.6 ;
        RECT 15.376 0 15.516 6.6 ;
        RECT 14.856 0 14.996 6.6 ;
        RECT 14.336 0 14.476 6.6 ;
        RECT 13.816 0 13.956 6.6 ;
        RECT 13.296 0 13.436 6.6 ;
        RECT 12.776 0 12.916 6.6 ;
        RECT 12.256 0 12.396 6.6 ;
        RECT 11.736 0 11.876 6.6 ;
        RECT 11.216 0 11.356 6.6 ;
        RECT 10.696 0 10.836 6.6 ;
        RECT 10.176 0 10.316 6.6 ;
        RECT 9.656 0 9.796 6.6 ;
        RECT 9.136 0 9.276 6.6 ;
        RECT 8.616 0 8.756 6.6 ;
        RECT 8.096 0 8.236 6.6 ;
        RECT 7.576 0 7.716 6.6 ;
        RECT 7.056 0 7.196 6.6 ;
        RECT 6.536 0 6.676 6.6 ;
        RECT 6.016 0 6.156 6.6 ;
        RECT 5.496 0 5.636 6.6 ;
        RECT 4.976 0 5.116 6.6 ;
        RECT 4.456 0 4.596 6.6 ;
        RECT 3.936 0 4.076 6.6 ;
        RECT 3.416 0 3.556 6.6 ;
        RECT 2.896 0 3.036 6.6 ;
        RECT 2.376 0 2.516 6.6 ;
        RECT 1.856 0 1.996 6.6 ;
        RECT 1.336 0 1.476 6.6 ;
    END
  END VSS
  PIN EN_N_CS_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 9.464286 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.956 0 24.096 6.6 ;
    END
  END EN_N_CS_I
  PIN CLK_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16192 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 22.916 0 23.056 6.6 ;
    END
  END CLK_O
  PIN EN_N_CR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 6.446429 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.696 0 23.836 6.6 ;
    END
  END EN_N_CR_I
  OBS
    LAYER CA ;
      RECT 0 0 25.172 6.6 ;
    LAYER M1 ;
      RECT 0 0 25.172 6.6 ;
    LAYER V1 ;
      RECT 0 0 25.172 6.6 ;
    LAYER M2 ;
      RECT 0 0 25.172 6.6 ;
    LAYER CB ;
      RECT 0 0 25.172 6.6 ;
    LAYER AY ;
      RECT 0 0 25.172 6.6 ;
    LAYER C1 ;
      RECT 18.236 0 18.376 6.6 ;
      RECT 18.235 1.82 18.376 1.9 ;
      RECT 24.996 0 25.136 6.6 ;
      RECT 24.736 0 24.876 6.6 ;
      RECT 24.476 0 24.616 6.6 ;
      RECT 24.216 0 24.356 6.6 ;
      RECT 23.956 0 24.096 6.6 ;
      RECT 23.696 0 23.836 6.6 ;
      RECT 23.436 0 23.576 0.72 ;
      RECT 23.436 0.84 23.576 5.04 ;
      RECT 23.436 5.16 23.576 6.6 ;
      RECT 23.176 0 23.316 6.6 ;
      RECT 22.916 0 23.056 6.6 ;
      RECT 22.656 0 22.796 6.6 ;
      RECT 22.396 0 22.536 0.72 ;
      RECT 22.396 0.84 22.536 2.16 ;
      RECT 22.396 2.28 22.536 5.04 ;
      RECT 22.396 5.16 22.536 6.6 ;
      RECT 22.136 0 22.276 6.6 ;
      RECT 21.876 0 22.016 0.72 ;
      RECT 21.876 0.84 22.016 2.16 ;
      RECT 21.876 2.28 22.016 5.76 ;
      RECT 21.876 5.88 22.016 6.6 ;
      RECT 21.616 0 21.756 6.6 ;
      RECT 21.356 0 21.496 6.6 ;
      RECT 21.096 0 21.236 6.6 ;
      RECT 20.836 0 20.976 2.16 ;
      RECT 20.836 2.28 20.976 2.62 ;
      RECT 20.836 2.7 20.976 5.04 ;
      RECT 20.836 5.16 20.976 6.6 ;
      RECT 20.576 0 20.716 6.6 ;
      RECT 20.316 0 20.456 6.6 ;
      RECT 20.056 0 20.196 6.6 ;
      RECT 19.796 0 19.936 6.6 ;
      RECT 19.536 0 19.676 6.6 ;
      RECT 19.276 0 19.416 6.6 ;
      RECT 19.016 0 19.156 6.6 ;
      RECT 18.756 0 18.896 6.6 ;
      RECT 18.496 0 18.636 6.6 ;
      RECT 17.976 0 18.116 6.6 ;
      RECT 17.716 0 17.856 6.6 ;
      RECT 17.456 0 17.596 6.6 ;
      RECT 17.196 0 17.336 6.6 ;
      RECT 16.936 0 17.076 6.6 ;
      RECT 16.676 0 16.816 6.6 ;
      RECT 16.416 0 16.556 6.6 ;
      RECT 16.156 0 16.296 6.6 ;
      RECT 15.896 0 16.036 6.6 ;
      RECT 15.636 0 15.776 6.6 ;
      RECT 15.376 0 15.516 6.6 ;
      RECT 15.116 0 15.256 6.6 ;
      RECT 14.856 0 14.996 6.6 ;
      RECT 14.596 0 14.736 6.6 ;
      RECT 14.336 0 14.476 6.6 ;
      RECT 14.076 0 14.216 6.6 ;
      RECT 13.816 0 13.956 6.6 ;
      RECT 13.556 0 13.696 6.6 ;
      RECT 13.296 0 13.436 6.6 ;
      RECT 13.036 0 13.176 6.6 ;
      RECT 12.776 0 12.916 6.6 ;
      RECT 12.516 0 12.656 6.6 ;
      RECT 12.256 0 12.396 6.6 ;
      RECT 11.996 0 12.136 6.6 ;
      RECT 11.736 0 11.876 6.6 ;
      RECT 11.476 0 11.616 6.6 ;
      RECT 11.216 0 11.356 6.6 ;
      RECT 10.956 0 11.096 6.6 ;
      RECT 10.696 0 10.836 6.6 ;
      RECT 10.436 0 10.576 6.6 ;
      RECT 10.176 0 10.316 6.6 ;
      RECT 9.916 0 10.056 6.6 ;
      RECT 9.656 0 9.796 6.6 ;
      RECT 9.396 0 9.536 6.6 ;
      RECT 9.136 0 9.276 6.6 ;
      RECT 8.876 0 9.016 6.6 ;
      RECT 8.616 0 8.756 6.6 ;
      RECT 8.356 0 8.496 0.72 ;
      RECT 8.356 0.84 8.496 1.44 ;
      RECT 8.356 1.56 8.496 6.6 ;
      RECT 8.096 0 8.236 6.6 ;
      RECT 7.836 0 7.976 6.6 ;
      RECT 7.576 0 7.716 6.6 ;
      RECT 7.316 0 7.456 6.6 ;
      RECT 7.056 0 7.196 6.6 ;
      RECT 6.796 0 6.936 6.6 ;
      RECT 6.536 0 6.676 6.6 ;
      RECT 6.276 0 6.416 0.72 ;
      RECT 6.276 0.84 6.416 5.04 ;
      RECT 6.276 5.16 6.416 6.6 ;
      RECT 6.016 0 6.156 6.6 ;
      RECT 5.756 0 5.896 6.6 ;
      RECT 5.496 0 5.636 6.6 ;
      RECT 5.236 0 5.376 6.6 ;
      RECT 4.976 0 5.116 6.6 ;
      RECT 4.716 0 4.856 6.6 ;
      RECT 4.456 0 4.596 6.6 ;
      RECT 4.196 0 4.336 6.6 ;
      RECT 3.936 0 4.076 6.6 ;
      RECT 3.676 0 3.816 6.6 ;
      RECT 3.416 0 3.556 6.6 ;
      RECT 3.156 0 3.296 1.44 ;
      RECT 3.156 1.56 3.296 2.88 ;
      RECT 3.156 3 3.296 4.32 ;
      RECT 3.156 4.44 3.296 6.6 ;
      RECT 2.896 0 3.036 6.6 ;
      RECT 2.636 0 2.776 0.72 ;
      RECT 2.636 0.84 2.776 4.32 ;
      RECT 2.636 4.44 2.776 5.76 ;
      RECT 2.636 5.88 2.776 6.6 ;
      RECT 2.376 0 2.516 6.6 ;
      RECT 2.116 0 2.256 6.6 ;
      RECT 1.856 0 1.996 6.6 ;
      RECT 1.596 0 1.736 6.6 ;
      RECT 1.336 0 1.476 6.6 ;
      RECT 1.076 0 1.216 1.44 ;
      RECT 1.076 1.56 1.216 2.88 ;
      RECT 1.076 4.44 1.216 6.6 ;
      RECT 0.816 0 0.956 6.6 ;
      RECT 0.556 0 0.696 6.6 ;
      RECT 0.296 0 0.436 6.6 ;
      RECT 0.036 0 0.176 6.6 ;
  END
END RIIO_RVT36G1_RESETGEN27

END LIBRARY
