VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


MACRO RIIO_EG1D80V_HPLVDS_RX_SLVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_HPLVDS_RX_SLVT28_V 0 0 ;
  SIZE 180 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN RTERM_TRIM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.348214 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.35 79.84 39.51 80 ;
    END
  END RTERM_TRIM_I[3]
  PIN RTERM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.401664 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 27.91 79.84 28.07 80 ;
    END
  END RTERM_EN_I
  PIN RTERM_TRIM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.419643 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 28.43 79.84 28.59 80 ;
    END
  END RTERM_TRIM_I[0]
  PIN RX_GAIN_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0944 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.184 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 386.518889 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 87.45 79.84 87.61 80 ;
    END
  END RX_GAIN_I[2]
  PIN EI_DETECT_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.01654 LAYER C1 ;
    ANTENNADIFFAREA 0.081 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 110.33 79.84 110.49 80 ;
    END
  END EI_DETECT_O
  PIN RX_CTLE_RES_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7585 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0416 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 690.423232 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 90.31 79.84 90.47 80 ;
    END
  END RX_CTLE_RES_I[1]
  PIN RX_CTLE_CAP_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7585 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0416 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 896.394949 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 89.53 79.84 89.69 80 ;
    END
  END RX_CTLE_CAP_I[3]
  PIN RX_CTLE_CAP_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7795 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0336 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.256 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 872.669697 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 89.01 79.84 89.17 80 ;
    END
  END RX_CTLE_CAP_I[2]
  PIN RX_CTLE_RES_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8215 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.208 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 687.192929 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 91.87 79.84 92.03 80 ;
    END
  END RX_CTLE_RES_I[4]
  PIN RX_CTLE_RES_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8005 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0496 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.232 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 688.269697 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 91.35 79.84 91.51 80 ;
    END
  END RX_CTLE_RES_I[3]
  PIN RX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8845 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1392 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 384.76 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 86.41 79.84 86.57 80 ;
    END
  END RX_EN_I
  PIN RX_CTLE_RES_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7795 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.02744 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.256 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 689.346465 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 90.83 79.84 90.99 80 ;
    END
  END RX_CTLE_RES_I[2]
  PIN RTERM_TRIM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.741071 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 32.07 79.84 32.23 80 ;
    END
  END RTERM_TRIM_I[1]
  PIN RX_CTLE_CAP_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8005 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0496 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.232 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 873.912121 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 88.49 79.84 88.65 80 ;
    END
  END RX_CTLE_CAP_I[1]
  PIN RTERM_TRIM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.544643 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.71 79.84 35.87 80 ;
    END
  END RTERM_TRIM_I[2]
  PIN RX_CTLE_RES_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8845 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1392 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 683.977778 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 93.43 79.84 93.59 80 ;
    END
  END RX_CTLE_RES_I[7]
  PIN A_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3851.735 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 4615.621 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 3859.61 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 2934.7608 LAYER JA ;
    ANTENNAPARTIALMETALAREA 4372.8408 LAYER QA ;
    ANTENNAPARTIALMETALAREA 3812.2008 LAYER QB ;
    ANTENNAPARTIALMETALAREA 1632.21795 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 76.332608 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 64.360384 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 165.568536 LAYER YS ;
    ANTENNAPARTIALCUTAREA 241.92 LAYER JV ;
    ANTENNAPARTIALCUTAREA 293.76 LAYER JW ;
    ANTENNAPARTIALCUTAREA 32.946144 LAYER A2 ;
    ANTENNADIFFAREA 889.8282 LAYER C4 ;
    ANTENNADIFFAREA 889.8282 LAYER C3 ;
    ANTENNADIFFAREA 889.8282 LAYER C5 ;
    ANTENNADIFFAREA 889.8282 LAYER JA ;
    ANTENNADIFFAREA 889.8282 LAYER QA ;
    ANTENNADIFFAREA 889.8282 LAYER QB ;
    ANTENNADIFFAREA 551.0762 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 2 24 87.6 28.8 ;
        RECT 81.4 0 86.2 2.4 ;
        RECT 75.2 0 80 2.4 ;
        RECT 69 0 73.8 2.4 ;
        RECT 62.8 0 67.6 2.4 ;
        RECT 56.6 0 61.4 2.4 ;
        RECT 50.4 0 55.2 2.4 ;
        RECT 44.2 0 49 2.4 ;
        RECT 38 0 42.8 2.4 ;
        RECT 31.8 0 36.6 2.4 ;
        RECT 25.6 0 30.4 2.4 ;
        RECT 19.4 0 24.2 2.4 ;
        RECT 13.2 0 18 2.4 ;
        RECT 7 0 11.8 2.4 ;
        RECT 0.8 0 5.6 2.4 ;
      LAYER QA ;
        RECT 81.4 0 86.2 2.4 ;
        RECT 75.2 0 80 2.4 ;
        RECT 69 0 73.8 2.4 ;
        RECT 62.8 0 67.6 2.4 ;
        RECT 56.6 0 61.4 2.4 ;
        RECT 50.4 0 55.2 2.4 ;
        RECT 44.2 0 49 2.4 ;
        RECT 38 0 42.8 2.4 ;
        RECT 31.8 0 36.6 2.4 ;
        RECT 25.6 0 30.4 2.4 ;
        RECT 19.4 0 24.2 2.4 ;
        RECT 13.2 0 18 2.4 ;
        RECT 7 0 11.8 2.4 ;
        RECT 0.8 0 5.6 2.4 ;
      LAYER JA ;
        RECT 81.4 0 86.2 2.4 ;
        RECT 75.2 0 80 2.4 ;
        RECT 69 0 73.8 2.4 ;
        RECT 62.8 0 67.6 2.4 ;
        RECT 56.6 0 61.4 2.4 ;
        RECT 50.4 0 55.2 2.4 ;
        RECT 44.2 0 49 2.4 ;
        RECT 38 0 42.8 2.4 ;
        RECT 31.8 0 36.6 2.4 ;
        RECT 25.6 0 30.4 2.4 ;
        RECT 19.4 0 24.2 2.4 ;
        RECT 13.2 0 18 2.4 ;
        RECT 7 0 11.8 2.4 ;
        RECT 0.8 0 5.6 2.4 ;
      LAYER C5 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
      LAYER C4 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
      LAYER C2 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 1.25 0 4.85 1.85 ;
      LAYER C3 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
    END
  END A_PAD_B
  PIN RX_CTLE_RES_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8635 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1168 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 685.039394 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 92.91 79.84 93.07 80 ;
    END
  END RX_CTLE_RES_I[6]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 0.8 75.2 5.6 80 ;
      LAYER QA ;
        RECT 0.8 75.2 5.6 80 ;
      LAYER JA ;
        RECT 0.8 75.2 5.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 13.2 75.2 18 80 ;
      LAYER QA ;
        RECT 13.2 75.2 18 80 ;
      LAYER JA ;
        RECT 13.2 75.2 18 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 25.6 75.2 30.4 80 ;
      LAYER QA ;
        RECT 25.6 75.2 30.4 80 ;
      LAYER JA ;
        RECT 25.6 75.2 30.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 38 75.2 42.8 80 ;
      LAYER QA ;
        RECT 38 75.2 42.8 80 ;
      LAYER JA ;
        RECT 38 75.2 42.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 50.4 75.2 55.2 80 ;
      LAYER QA ;
        RECT 50.4 75.2 55.2 80 ;
      LAYER JA ;
        RECT 50.4 75.2 55.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 62.8 75.2 67.6 80 ;
      LAYER QA ;
        RECT 62.8 75.2 67.6 80 ;
      LAYER JA ;
        RECT 62.8 75.2 67.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 75.2 80 80 ;
      LAYER QA ;
        RECT 75.2 75.2 80 80 ;
      LAYER JA ;
        RECT 75.2 75.2 80 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 87.6 75.2 92.4 80 ;
      LAYER QA ;
        RECT 87.6 75.2 92.4 80 ;
      LAYER JA ;
        RECT 87.6 75.2 92.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 100 75.2 104.8 80 ;
      LAYER QA ;
        RECT 100 75.2 104.8 80 ;
      LAYER JA ;
        RECT 100 75.2 104.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 112.4 75.2 117.2 80 ;
      LAYER QA ;
        RECT 112.4 75.2 117.2 80 ;
      LAYER JA ;
        RECT 112.4 75.2 117.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 124.8 75.2 129.6 80 ;
      LAYER QA ;
        RECT 124.8 75.2 129.6 80 ;
      LAYER JA ;
        RECT 124.8 75.2 129.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 137.2 75.2 142 80 ;
      LAYER QA ;
        RECT 137.2 75.2 142 80 ;
      LAYER JA ;
        RECT 137.2 75.2 142 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 149.6 75.2 154.4 80 ;
      LAYER QA ;
        RECT 149.6 75.2 154.4 80 ;
      LAYER JA ;
        RECT 149.6 75.2 154.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 162 75.2 166.8 80 ;
      LAYER QA ;
        RECT 162 75.2 166.8 80 ;
      LAYER JA ;
        RECT 162 75.2 166.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 174.4 75.2 179.2 80 ;
      LAYER QA ;
        RECT 174.4 75.2 179.2 80 ;
      LAYER JA ;
        RECT 174.4 75.2 179.2 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 67.4 180 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 180 53.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 7 75.2 11.8 80 ;
      LAYER QA ;
        RECT 7 75.2 11.8 80 ;
      LAYER JA ;
        RECT 7 75.2 11.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 19.4 75.2 24.2 80 ;
      LAYER QA ;
        RECT 19.4 75.2 24.2 80 ;
      LAYER JA ;
        RECT 19.4 75.2 24.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 31.8 75.2 36.6 80 ;
      LAYER QA ;
        RECT 31.8 75.2 36.6 80 ;
      LAYER JA ;
        RECT 31.8 75.2 36.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 44.2 75.2 49 80 ;
      LAYER QA ;
        RECT 44.2 75.2 49 80 ;
      LAYER JA ;
        RECT 44.2 75.2 49 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 56.6 75.2 61.4 80 ;
      LAYER QA ;
        RECT 56.6 75.2 61.4 80 ;
      LAYER JA ;
        RECT 56.6 75.2 61.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 69 75.2 73.8 80 ;
      LAYER QA ;
        RECT 69 75.2 73.8 80 ;
      LAYER JA ;
        RECT 69 75.2 73.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 81.4 75.2 86.2 80 ;
      LAYER QA ;
        RECT 81.4 75.2 86.2 80 ;
      LAYER JA ;
        RECT 81.4 75.2 86.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 93.8 75.2 98.6 80 ;
      LAYER QA ;
        RECT 93.8 75.2 98.6 80 ;
      LAYER JA ;
        RECT 93.8 75.2 98.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 106.2 75.2 111 80 ;
      LAYER QA ;
        RECT 106.2 75.2 111 80 ;
      LAYER JA ;
        RECT 106.2 75.2 111 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 118.6 75.2 123.4 80 ;
      LAYER QA ;
        RECT 118.6 75.2 123.4 80 ;
      LAYER JA ;
        RECT 118.6 75.2 123.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 131 75.2 135.8 80 ;
      LAYER QA ;
        RECT 131 75.2 135.8 80 ;
      LAYER JA ;
        RECT 131 75.2 135.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 143.4 75.2 148.2 80 ;
      LAYER QA ;
        RECT 143.4 75.2 148.2 80 ;
      LAYER JA ;
        RECT 143.4 75.2 148.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 155.8 75.2 160.6 80 ;
      LAYER QA ;
        RECT 155.8 75.2 160.6 80 ;
      LAYER JA ;
        RECT 155.8 75.2 160.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 168.2 75.2 173 80 ;
      LAYER QA ;
        RECT 168.2 75.2 173 80 ;
      LAYER JA ;
        RECT 168.2 75.2 173 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 61.2 180 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 180 59.8 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 180 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 180 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 180 10.2 ;
    END
  END VSSIO
  PIN B_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2385.0375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1287.3555 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 2651.475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 2325.6408 LAYER JA ;
    ANTENNAPARTIALMETALAREA 3087.8808 LAYER QA ;
    ANTENNAPARTIALMETALAREA 3196.3608 LAYER QB ;
    ANTENNAPARTIALMETALAREA 35.36175 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 24.45168 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.602784 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 132.146316 LAYER YS ;
    ANTENNAPARTIALCUTAREA 172.8 LAYER JV ;
    ANTENNAPARTIALCUTAREA 224.64 LAYER JW ;
    ANTENNAPARTIALCUTAREA 10.82224 LAYER A2 ;
    ANTENNADIFFAREA 721.7962 LAYER C4 ;
    ANTENNADIFFAREA 334.12 LAYER C3 ;
    ANTENNADIFFAREA 721.7962 LAYER C5 ;
    ANTENNADIFFAREA 721.7962 LAYER JA ;
    ANTENNADIFFAREA 721.7962 LAYER QA ;
    ANTENNADIFFAREA 721.7962 LAYER QB ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 174.417 0 179.217 2.4 ;
        RECT 92.4 24 178 28.8 ;
        RECT 168.217 0 173.017 2.4 ;
        RECT 162.017 0 166.817 2.4 ;
        RECT 155.817 0 160.617 2.4 ;
        RECT 149.617 0 154.417 2.4 ;
        RECT 143.417 0 148.217 2.4 ;
        RECT 137.217 0 142.017 2.4 ;
        RECT 131.017 0 135.817 2.4 ;
        RECT 124.817 0 129.617 2.4 ;
        RECT 118.617 0 123.417 2.4 ;
        RECT 112.417 0 117.217 2.4 ;
        RECT 106.217 0 111.017 2.4 ;
        RECT 100.017 0 104.817 2.4 ;
        RECT 93.817 0 98.617 2.4 ;
      LAYER QA ;
        RECT 174.417 0 179.217 2.4 ;
        RECT 168.217 0 173.017 2.4 ;
        RECT 162.017 0 166.817 2.4 ;
        RECT 155.817 0 160.617 2.4 ;
        RECT 149.617 0 154.417 2.4 ;
        RECT 143.417 0 148.217 2.4 ;
        RECT 137.217 0 142.017 2.4 ;
        RECT 131.017 0 135.817 2.4 ;
        RECT 124.817 0 129.617 2.4 ;
        RECT 118.617 0 123.417 2.4 ;
        RECT 112.417 0 117.217 2.4 ;
        RECT 106.217 0 111.017 2.4 ;
        RECT 100.017 0 104.817 2.4 ;
        RECT 93.817 0 98.617 2.4 ;
      LAYER JA ;
        RECT 174.417 0 179.217 2.4 ;
        RECT 168.217 0 173.017 2.4 ;
        RECT 162.017 0 166.817 2.4 ;
        RECT 155.817 0 160.617 2.4 ;
        RECT 149.617 0 154.417 2.4 ;
        RECT 143.417 0 148.217 2.4 ;
        RECT 137.217 0 142.017 2.4 ;
        RECT 131.017 0 135.817 2.4 ;
        RECT 124.817 0 129.617 2.4 ;
        RECT 118.617 0 123.417 2.4 ;
        RECT 112.417 0 117.217 2.4 ;
        RECT 106.217 0 111.017 2.4 ;
        RECT 100.017 0 104.817 2.4 ;
        RECT 93.817 0 98.617 2.4 ;
      LAYER C5 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C4 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C2 ;
        RECT 175.15 0 178.75 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C3 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
    END
  END B_PAD_B
  PIN EI_DETECT_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 67.95 79.84 68.11 80 ;
    END
  END EI_DETECT_EN_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 180 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 180 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 180 16.4 ;
    END
  END VDDIO
  PIN DI_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNADIFFAREA 0.16192 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 67.43 79.84 67.59 80 ;
    END
  END DI_O
  PIN RX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 64.31 79.84 64.47 80 ;
    END
  END RX_VCM_EN_I
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.408 LAYER C4 ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER C4 ;
        RECT 0 39.575 180 40.825 ;
    END
  END VBIAS
  PIN RX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C1 ;
      ANTENNAMAXAREACAR 11.598214 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 69.51 79.84 69.67 80 ;
    END
  END RX_POL_I
  PIN RX_GAIN_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8215 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.208 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 385.255556 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 87.97 79.84 88.13 80 ;
    END
  END RX_GAIN_I[3]
  PIN RX_CTLE_RES_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0944 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.184 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 686.116162 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 92.39 79.84 92.55 80 ;
    END
  END RX_CTLE_RES_I[5]
  PIN RX_GAIN_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8635 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1168 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 385.923333 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 86.93 79.84 87.09 80 ;
    END
  END RX_GAIN_I[1]
  OBS
    LAYER CA ;
      RECT 0 0 180 80 ;
    LAYER M1 ;
      RECT 0 0 180 80 ;
    LAYER V1 ;
      RECT 0 0 180 80 ;
    LAYER M2 ;
      RECT 0 0 180 80 ;
    LAYER A1 ;
      RECT 0 0 180 80 ;
    LAYER C2 ;
      RECT 0 0 180 80 ;
    LAYER CB ;
      RECT 0 0 180 80 ;
    LAYER JV ;
      RECT 0 0 180 80 ;
    LAYER YS ;
      RECT 0 0 180 80 ;
    LAYER JW ;
      RECT 0 0 180 80 ;
    LAYER QB ;
      RECT 0 0 180 80 ;
    LAYER QA ;
      RECT 0 0 180 80 ;
    LAYER JA ;
      RECT 0 0 180 80 ;
    LAYER AY ;
      RECT 0 0 180 80 ;
    LAYER C1 ;
      RECT 0 0 180 80 ;
    LAYER C5 ;
      RECT 0 0 180 80 ;
    LAYER C4 ;
      RECT 0 0 180 80 ;
    LAYER C3 ;
      RECT 0 0 180 80 ;
    LAYER A4 ;
      RECT 0 0 180 80 ;
    LAYER A3 ;
      RECT 0 0 180 80 ;
    LAYER A2 ;
      RECT 0 0 180 80 ;
  END
END RIIO_EG1D80V_HPLVDS_RX_SLVT28_V

MACRO RIIO_EG1D80V_HPLVDS_TX_SLVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_HPLVDS_TX_SLVT28_V 0 0 ;
  SIZE 180 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN TX_FFE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02128 LAYER C1 ;
      ANTENNAMAXAREACAR 14.671992 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 49.23 79.84 49.39 80 ;
    END
  END TX_FFE_I
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.408 LAYER C4 ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER C4 ;
        RECT 0 39.575 180 40.825 ;
    END
  END VBIAS
  PIN RTERM_TRIM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.348214 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.35 79.84 39.51 80 ;
    END
  END RTERM_TRIM_I[3]
  PIN RTERM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.401664 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 27.91 79.84 28.07 80 ;
    END
  END RTERM_EN_I
  PIN RTERM_TRIM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.419643 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 28.43 79.84 28.59 80 ;
    END
  END RTERM_TRIM_I[0]
  PIN TX_BIAS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.517857 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 18.03 79.84 18.19 80 ;
    END
  END TX_BIAS_I[0]
  PIN RX_GAIN_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0944 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.184 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 386.518889 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 87.45 79.84 87.61 80 ;
    END
  END RX_GAIN_I[2]
  PIN TX_EI_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0112 LAYER C1 ;
      ANTENNAMAXAREACAR 22.714286 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 45.33 79.84 45.49 80 ;
    END
  END TX_EI_I
  PIN EI_DETECT_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.01654 LAYER C1 ;
    ANTENNADIFFAREA 0.081 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 110.33 79.84 110.49 80 ;
    END
  END EI_DETECT_O
  PIN RX_CTLE_RES_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7585 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0416 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 690.423232 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 90.31 79.84 90.47 80 ;
    END
  END RX_CTLE_RES_I[1]
  PIN RX_CTLE_CAP_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7585 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0416 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 896.394949 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 89.53 79.84 89.69 80 ;
    END
  END RX_CTLE_CAP_I[3]
  PIN RX_CTLE_CAP_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7795 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0336 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.256 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 872.669697 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 89.01 79.84 89.17 80 ;
    END
  END RX_CTLE_CAP_I[2]
  PIN TX_VCM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.446429 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 48.19 79.84 48.35 80 ;
    END
  END TX_VCM_I[3]
  PIN RX_CTLE_RES_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8215 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.208 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 687.192929 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 91.87 79.84 92.03 80 ;
    END
  END RX_CTLE_RES_I[4]
  PIN RX_CTLE_RES_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8005 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0496 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.232 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 688.269697 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 91.35 79.84 91.51 80 ;
    END
  END RX_CTLE_RES_I[3]
  PIN RX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8845 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1392 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 384.76 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 86.41 79.84 86.57 80 ;
    END
  END RX_EN_I
  PIN RX_CTLE_RES_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7795 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.02744 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.256 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 689.346465 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 90.83 79.84 90.99 80 ;
    END
  END RX_CTLE_RES_I[2]
  PIN TX_VCM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.517857 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 59.11 79.84 59.27 80 ;
    END
  END TX_VCM_I[0]
  PIN TX_BIAS_OD_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.23 79.84 23.39 80 ;
    END
  END TX_BIAS_OD_I
  PIN RTERM_TRIM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.741071 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 32.07 79.84 32.23 80 ;
    END
  END RTERM_TRIM_I[1]
  PIN RX_CTLE_CAP_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8005 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0496 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.232 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 873.912121 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 88.49 79.84 88.65 80 ;
    END
  END RX_CTLE_CAP_I[1]
  PIN TX_BIAS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.839286 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.39 79.84 14.55 80 ;
    END
  END TX_BIAS_I[1]
  PIN TX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.304261 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.59 79.84 19.75 80 ;
    END
  END TX_EN_I
  PIN TX_BIAS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.642857 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.75 79.84 10.91 80 ;
    END
  END TX_BIAS_I[2]
  PIN TX_BIAS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.446429 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 7.11 79.84 7.27 80 ;
    END
  END TX_BIAS_I[3]
  PIN RTERM_TRIM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.544643 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.71 79.84 35.87 80 ;
    END
  END RTERM_TRIM_I[2]
  PIN RX_CTLE_RES_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8845 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1392 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 683.977778 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 93.43 79.84 93.59 80 ;
    END
  END RX_CTLE_RES_I[7]
  PIN A_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3851.735 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 4615.621 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 3859.61 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 2934.7608 LAYER JA ;
    ANTENNAPARTIALMETALAREA 4372.8408 LAYER QA ;
    ANTENNAPARTIALMETALAREA 3812.2008 LAYER QB ;
    ANTENNAPARTIALMETALAREA 1632.21795 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 76.332608 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 64.360384 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 165.568536 LAYER YS ;
    ANTENNAPARTIALCUTAREA 241.92 LAYER JV ;
    ANTENNAPARTIALCUTAREA 293.76 LAYER JW ;
    ANTENNAPARTIALCUTAREA 32.946144 LAYER A2 ;
    ANTENNADIFFAREA 997.3482 LAYER C4 ;
    ANTENNADIFFAREA 997.3482 LAYER C3 ;
    ANTENNADIFFAREA 997.3482 LAYER C5 ;
    ANTENNADIFFAREA 997.3482 LAYER JA ;
    ANTENNADIFFAREA 997.3482 LAYER QA ;
    ANTENNADIFFAREA 997.3482 LAYER QB ;
    ANTENNADIFFAREA 551.0762 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 2 24 87.6 28.8 ;
        RECT 81.4 0 86.2 2.4 ;
        RECT 75.2 0 80 2.4 ;
        RECT 69 0 73.8 2.4 ;
        RECT 62.8 0 67.6 2.4 ;
        RECT 56.6 0 61.4 2.4 ;
        RECT 50.4 0 55.2 2.4 ;
        RECT 44.2 0 49 2.4 ;
        RECT 38 0 42.8 2.4 ;
        RECT 31.8 0 36.6 2.4 ;
        RECT 25.6 0 30.4 2.4 ;
        RECT 19.4 0 24.2 2.4 ;
        RECT 13.2 0 18 2.4 ;
        RECT 7 0 11.8 2.4 ;
        RECT 0.8 0 5.6 2.4 ;
      LAYER QA ;
        RECT 81.4 0 86.2 2.4 ;
        RECT 75.2 0 80 2.4 ;
        RECT 69 0 73.8 2.4 ;
        RECT 62.8 0 67.6 2.4 ;
        RECT 56.6 0 61.4 2.4 ;
        RECT 50.4 0 55.2 2.4 ;
        RECT 44.2 0 49 2.4 ;
        RECT 38 0 42.8 2.4 ;
        RECT 31.8 0 36.6 2.4 ;
        RECT 25.6 0 30.4 2.4 ;
        RECT 19.4 0 24.2 2.4 ;
        RECT 13.2 0 18 2.4 ;
        RECT 7 0 11.8 2.4 ;
        RECT 0.8 0 5.6 2.4 ;
      LAYER JA ;
        RECT 81.4 0 86.2 2.4 ;
        RECT 75.2 0 80 2.4 ;
        RECT 69 0 73.8 2.4 ;
        RECT 62.8 0 67.6 2.4 ;
        RECT 56.6 0 61.4 2.4 ;
        RECT 50.4 0 55.2 2.4 ;
        RECT 44.2 0 49 2.4 ;
        RECT 38 0 42.8 2.4 ;
        RECT 31.8 0 36.6 2.4 ;
        RECT 25.6 0 30.4 2.4 ;
        RECT 19.4 0 24.2 2.4 ;
        RECT 13.2 0 18 2.4 ;
        RECT 7 0 11.8 2.4 ;
        RECT 0.8 0 5.6 2.4 ;
      LAYER C5 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
      LAYER C3 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
      LAYER C4 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
      LAYER C2 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 1.25 0 4.85 1.85 ;
    END
  END A_PAD_B
  PIN RX_CTLE_RES_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8635 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1168 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 685.039394 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 92.91 79.84 93.07 80 ;
    END
  END RX_CTLE_RES_I[6]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    ANTENNAPARTIALMETALAREA 2027.52 LAYER QB ;
    ANTENNAPARTIALMETALAREA 126.72 LAYER QA ;
    ANTENNAPARTIALCUTAREA 5.76 LAYER JV ;
    ANTENNAPARTIALCUTAREA 17.28 LAYER JW ;
    ANTENNADIFFAREA 59.00996 LAYER QA ;
    ANTENNADIFFAREA 59.00996 LAYER QB ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 8.91504 LAYER QA ;
      ANTENNAGATEAREA 8.91504 LAYER QB ;
      ANTENNAMAXAREACAR 28.928273 LAYER QA ;
      ANTENNAMAXAREACAR 45.082688 LAYER QB ;
      ANTENNAMAXCUTCAR 0.583938 LAYER JW ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 168.2 75.2 173 80 ;
        RECT 155.8 75.2 160.6 80 ;
        RECT 143.4 75.2 148.2 80 ;
        RECT 131 75.2 135.8 80 ;
        RECT 118.6 75.2 123.4 80 ;
        RECT 106.2 75.2 111 80 ;
        RECT 93.8 75.2 98.6 80 ;
        RECT 81.4 75.2 86.2 80 ;
        RECT 69 75.2 73.8 80 ;
        RECT 56.6 75.2 61.4 80 ;
        RECT 44.2 75.2 49 80 ;
        RECT 31.8 75.2 36.6 80 ;
        RECT 19.4 75.2 24.2 80 ;
        RECT 7 75.2 11.8 80 ;
      LAYER QA ;
        RECT 168.2 75.2 173 80 ;
        RECT 155.8 75.2 160.6 80 ;
        RECT 143.4 75.2 148.2 80 ;
        RECT 131 75.2 135.8 80 ;
        RECT 118.6 75.2 123.4 80 ;
        RECT 106.2 75.2 111 80 ;
        RECT 93.8 75.2 98.6 80 ;
        RECT 81.4 75.2 86.2 80 ;
        RECT 69 75.2 73.8 80 ;
        RECT 56.6 75.2 61.4 80 ;
        RECT 44.2 75.2 49 80 ;
        RECT 31.8 75.2 36.6 80 ;
        RECT 19.4 75.2 24.2 80 ;
        RECT 7 75.2 11.8 80 ;
      LAYER JA ;
        RECT 168.2 75.2 173 80 ;
        RECT 155.8 75.2 160.6 80 ;
        RECT 143.4 75.2 148.2 80 ;
        RECT 131 75.2 135.8 80 ;
        RECT 118.6 75.2 123.4 80 ;
        RECT 106.2 75.2 111 80 ;
        RECT 93.8 75.2 98.6 80 ;
        RECT 81.4 75.2 86.2 80 ;
        RECT 69 75.2 73.8 80 ;
        RECT 56.6 75.2 61.4 80 ;
        RECT 44.2 75.2 49 80 ;
        RECT 31.8 75.2 36.6 80 ;
        RECT 19.4 75.2 24.2 80 ;
        RECT 7 75.2 11.8 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 180 59.8 ;
        RECT 0 61.2 180 66 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    ANTENNAPARTIALMETALAREA 2050.56 LAYER QB ;
    ANTENNAPARTIALMETALAREA 126.72 LAYER QA ;
    ANTENNAPARTIALCUTAREA 5.76 LAYER JV ;
    ANTENNAPARTIALCUTAREA 17.28 LAYER JW ;
    ANTENNADIFFAREA 98.917132 LAYER QA ;
    ANTENNADIFFAREA 98.917132 LAYER QB ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.11104 LAYER QA ;
      ANTENNAGATEAREA 1.11104 LAYER QB ;
      ANTENNAMAXAREACAR 2.326083 LAYER QB ;
      ANTENNAMAXCUTCAR 0.276457 LAYER JW ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 174.4 75.2 179.2 80 ;
        RECT 162 75.2 166.8 80 ;
        RECT 149.6 75.2 154.4 80 ;
        RECT 137.2 75.2 142 80 ;
        RECT 124.8 75.2 129.6 80 ;
        RECT 112.4 75.2 117.2 80 ;
        RECT 100 75.2 104.8 80 ;
        RECT 87.6 75.2 92.4 80 ;
        RECT 75.2 75.2 80 80 ;
        RECT 62.8 75.2 67.6 80 ;
        RECT 50.4 75.2 55.2 80 ;
        RECT 38 75.2 42.8 80 ;
        RECT 25.6 75.2 30.4 80 ;
        RECT 13.2 75.2 18 80 ;
        RECT 0.8 75.2 5.6 80 ;
      LAYER QA ;
        RECT 174.4 75.2 179.2 80 ;
        RECT 162 75.2 166.8 80 ;
        RECT 149.6 75.2 154.4 80 ;
        RECT 137.2 75.2 142 80 ;
        RECT 124.8 75.2 129.6 80 ;
        RECT 112.4 75.2 117.2 80 ;
        RECT 100 75.2 104.8 80 ;
        RECT 87.6 75.2 92.4 80 ;
        RECT 75.2 75.2 80 80 ;
        RECT 62.8 75.2 67.6 80 ;
        RECT 50.4 75.2 55.2 80 ;
        RECT 38 75.2 42.8 80 ;
        RECT 25.6 75.2 30.4 80 ;
        RECT 13.2 75.2 18 80 ;
        RECT 0.8 75.2 5.6 80 ;
      LAYER JA ;
        RECT 174.4 75.2 179.2 80 ;
        RECT 162 75.2 166.8 80 ;
        RECT 149.6 75.2 154.4 80 ;
        RECT 137.2 75.2 142 80 ;
        RECT 124.8 75.2 129.6 80 ;
        RECT 112.4 75.2 117.2 80 ;
        RECT 100 75.2 104.8 80 ;
        RECT 87.6 75.2 92.4 80 ;
        RECT 75.2 75.2 80 80 ;
        RECT 62.8 75.2 67.6 80 ;
        RECT 50.4 75.2 55.2 80 ;
        RECT 38 75.2 42.8 80 ;
        RECT 25.6 75.2 30.4 80 ;
        RECT 13.2 75.2 18 80 ;
        RECT 0.8 75.2 5.6 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 180 53.6 ;
        RECT 0 67.4 180 72.2 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    ANTENNAPARTIALMETALAREA 1728 LAYER QB ;
    ANTENNADIFFAREA 574.7898 LAYER QB ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.048 LAYER QB ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 5.4 180 10.2 ;
        RECT 0 17.8 180 22.6 ;
        RECT 0 42.6 180 47.4 ;
    END
  END VSSIO
  PIN B_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2385.0375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1287.3555 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 2651.475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 2325.6408 LAYER JA ;
    ANTENNAPARTIALMETALAREA 3087.8808 LAYER QA ;
    ANTENNAPARTIALMETALAREA 3196.3608 LAYER QB ;
    ANTENNAPARTIALMETALAREA 35.36175 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 24.45168 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.602784 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 132.146316 LAYER YS ;
    ANTENNAPARTIALCUTAREA 172.8 LAYER JV ;
    ANTENNAPARTIALCUTAREA 224.64 LAYER JW ;
    ANTENNAPARTIALCUTAREA 10.82224 LAYER A2 ;
    ANTENNADIFFAREA 775.5562 LAYER C4 ;
    ANTENNADIFFAREA 387.88 LAYER C3 ;
    ANTENNADIFFAREA 775.5562 LAYER C5 ;
    ANTENNADIFFAREA 775.5562 LAYER JA ;
    ANTENNADIFFAREA 775.5562 LAYER QA ;
    ANTENNADIFFAREA 775.5562 LAYER QB ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 174.417 0 179.217 2.4 ;
        RECT 92.4 24 178 28.8 ;
        RECT 168.217 0 173.017 2.4 ;
        RECT 162.017 0 166.817 2.4 ;
        RECT 155.817 0 160.617 2.4 ;
        RECT 149.617 0 154.417 2.4 ;
        RECT 143.417 0 148.217 2.4 ;
        RECT 137.217 0 142.017 2.4 ;
        RECT 131.017 0 135.817 2.4 ;
        RECT 124.817 0 129.617 2.4 ;
        RECT 118.617 0 123.417 2.4 ;
        RECT 112.417 0 117.217 2.4 ;
        RECT 106.217 0 111.017 2.4 ;
        RECT 100.017 0 104.817 2.4 ;
        RECT 93.817 0 98.617 2.4 ;
      LAYER QA ;
        RECT 174.417 0 179.217 2.4 ;
        RECT 168.217 0 173.017 2.4 ;
        RECT 162.017 0 166.817 2.4 ;
        RECT 155.817 0 160.617 2.4 ;
        RECT 149.617 0 154.417 2.4 ;
        RECT 143.417 0 148.217 2.4 ;
        RECT 137.217 0 142.017 2.4 ;
        RECT 131.017 0 135.817 2.4 ;
        RECT 124.817 0 129.617 2.4 ;
        RECT 118.617 0 123.417 2.4 ;
        RECT 112.417 0 117.217 2.4 ;
        RECT 106.217 0 111.017 2.4 ;
        RECT 100.017 0 104.817 2.4 ;
        RECT 93.817 0 98.617 2.4 ;
      LAYER JA ;
        RECT 174.417 0 179.217 2.4 ;
        RECT 168.217 0 173.017 2.4 ;
        RECT 162.017 0 166.817 2.4 ;
        RECT 155.817 0 160.617 2.4 ;
        RECT 149.617 0 154.417 2.4 ;
        RECT 143.417 0 148.217 2.4 ;
        RECT 137.217 0 142.017 2.4 ;
        RECT 131.017 0 135.817 2.4 ;
        RECT 124.817 0 129.617 2.4 ;
        RECT 118.617 0 123.417 2.4 ;
        RECT 112.417 0 117.217 2.4 ;
        RECT 106.217 0 111.017 2.4 ;
        RECT 100.017 0 104.817 2.4 ;
        RECT 93.817 0 98.617 2.4 ;
      LAYER C5 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C3 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C4 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C2 ;
        RECT 175.15 0 178.75 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
    END
  END B_PAD_B
  PIN EI_DETECT_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 67.95 79.84 68.11 80 ;
    END
  END EI_DETECT_EN_I
  PIN TX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.304261 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 60.67 79.84 60.83 80 ;
    END
  END TX_VCM_EN_I
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C1 ;
      ANTENNAMAXAREACAR 11.288393 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.99 79.84 43.15 80 ;
    END
  END DO_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    ANTENNAPARTIALMETALAREA 1728 LAYER QB ;
    ANTENNADIFFAREA 553.7642 LAYER QB ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 11.6 180 16.4 ;
        RECT 0 30.2 180 35 ;
        RECT 0 36.4 180 41.2 ;
    END
  END VDDIO
  PIN DI_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNADIFFAREA 0.16192 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 67.43 79.84 67.59 80 ;
    END
  END DI_O
  PIN RX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 64.31 79.84 64.47 80 ;
    END
  END RX_VCM_EN_I
  PIN TX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C1 ;
      ANTENNAMAXAREACAR 12.119643 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.47 79.84 42.63 80 ;
    END
  END TX_POL_I
  PIN RX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C1 ;
      ANTENNAMAXAREACAR 11.598214 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 69.51 79.84 69.67 80 ;
    END
  END RX_POL_I
  PIN RX_GAIN_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8215 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.208 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 385.255556 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 87.97 79.84 88.13 80 ;
    END
  END RX_GAIN_I[3]
  PIN RX_CTLE_RES_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0944 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.184 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 686.116162 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 92.39 79.84 92.55 80 ;
    END
  END RX_CTLE_RES_I[5]
  PIN RX_GAIN_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8635 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1168 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 385.923333 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 86.93 79.84 87.09 80 ;
    END
  END RX_GAIN_I[1]
  PIN TX_VCM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.839286 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 55.47 79.84 55.63 80 ;
    END
  END TX_VCM_I[1]
  PIN TX_VCM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.642857 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 51.83 79.84 51.99 80 ;
    END
  END TX_VCM_I[2]
  OBS
    LAYER CA ;
      RECT 0 0 180 80 ;
    LAYER M1 ;
      RECT 0 0 180 80 ;
    LAYER V1 ;
      RECT 0 0 180 80 ;
    LAYER M2 ;
      RECT 0 0 180 80 ;
    LAYER A1 ;
      RECT 0 0 180 80 ;
    LAYER C2 ;
      RECT 0 0 180 80 ;
    LAYER CB ;
      RECT 0 0 180 80 ;
    LAYER JV ;
      RECT 0 0 180 80 ;
    LAYER YS ;
      RECT 0 0 180 80 ;
    LAYER JW ;
      RECT 0 0 180 80 ;
    LAYER QB ;
      RECT 0 0 180 80 ;
    LAYER QA ;
      RECT 0 0 180 80 ;
    LAYER JA ;
      RECT 0 0 180 80 ;
    LAYER AY ;
      RECT 0 0 180 80 ;
    LAYER C1 ;
      RECT 0 0 180 80 ;
    LAYER C5 ;
      RECT 0 0 180 80 ;
    LAYER C4 ;
      RECT 0 0 180 80 ;
    LAYER C3 ;
      RECT 0 0 180 80 ;
    LAYER A4 ;
      RECT 0 0 180 80 ;
    LAYER A3 ;
      RECT 0 0 180 80 ;
    LAYER A2 ;
      RECT 0 0 180 80 ;
  END
END RIIO_EG1D80V_HPLVDS_TX_SLVT28_V

MACRO RIIO_EG1D80V_RTERMCAL_HVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_HVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.564137 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.2 79.86 40.34 80 ;
    END
  END D_IOSG_I[10]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2212 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.36 79.86 5.5 80 ;
    END
  END RESULT_O[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.84 79.86 4.98 80 ;
    END
  END RESULT_O[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.336729 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.4 79.86 19.54 80 ;
    END
  END MODE_I[1]
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.869565 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.04 79.86 23.18 80 ;
    END
  END MODE_I[0]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.058036 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.92 79.86 7.06 80 ;
    END
  END D_LVDS_I[3]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.736607 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.56 79.86 10.7 80 ;
    END
  END D_LVDS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 68.1725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 493.9475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 364.8 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 235.02 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.5176 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JV ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JW ;
    ANTENNAPARTIALCUTAREA 7.031552 LAYER A2 ;
    ANTENNADIFFAREA 167.0608 LAYER C4 ;
    ANTENNADIFFAREA 167.0608 LAYER C3 ;
    ANTENNADIFFAREA 167.0608 LAYER C5 ;
    ANTENNADIFFAREA 167.0608 LAYER JA ;
    ANTENNADIFFAREA 167.0608 LAYER QA ;
    ANTENNADIFFAREA 167.0608 LAYER QB ;
    ANTENNADIFFAREA 167.0608 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
        RECT 2 24 58 28.8 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
    END
  END PAD_B
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.84 79.86 30.98 80 ;
    END
  END VDDQ
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.450893 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.2 79.86 14.34 80 ;
    END
  END D_LVDS_I[1]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.129464 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.84 79.86 17.98 80 ;
    END
  END D_LVDS_I[0]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.637946 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.68 79.86 39.82 80 ;
    END
  END D_IOSG_I[9]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.518659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.16 79.86 39.3 80 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.594022 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.64 79.86 38.78 80 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.369792 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.12 79.86 38.26 80 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.446458 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.6 79.86 37.74 80 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.136806 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.08 79.86 37.22 80 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.214583 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.56 79.86 36.7 80 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.670735 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.04 79.86 36.18 80 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.747794 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.52 79.86 35.66 80 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C1 ;
      ANTENNAMAXAREACAR 2.443131 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.8 79.86 42.94 80 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C1 ;
      ANTENNAMAXAREACAR 2.582738 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.28 79.86 42.42 80 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C1 ;
      ANTENNAMAXAREACAR 2.733211 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.76 79.86 41.9 80 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.179861 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.24 79.86 41.38 80 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.253194 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.72 79.86 40.86 80 ;
    END
  END D_IOSG_I[11]
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.32 79.86 30.46 80 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_RTERMCAL_HVT28_V

MACRO RIIO_EG1D80V_RTERMCAL_LLHVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_LLHVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.564137 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.2 79.86 40.34 80 ;
    END
  END D_IOSG_I[10]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2212 LAYER C1 ;
    ANTENNADIFFAREA 0.03864 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.36 79.86 5.5 80 ;
    END
  END RESULT_O[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNADIFFAREA 0.03864 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.84 79.86 4.98 80 ;
    END
  END RESULT_O[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.044 LAYER C1 ;
      ANTENNAMAXAREACAR 22.719659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.4 79.86 19.54 80 ;
    END
  END MODE_I[1]
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0184 LAYER C1 ;
      ANTENNAMAXAREACAR 19.954348 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.04 79.86 23.18 80 ;
    END
  END MODE_I[0]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C1 ;
      ANTENNAMAXAREACAR 59.65625 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.92 79.86 7.06 80 ;
    END
  END D_LVDS_I[3]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C1 ;
      ANTENNAMAXAREACAR 59.65625 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.56 79.86 10.7 80 ;
    END
  END D_LVDS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 68.1725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 493.9475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 364.8 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 235.02 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.5176 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JV ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JW ;
    ANTENNAPARTIALCUTAREA 7.031552 LAYER A2 ;
    ANTENNADIFFAREA 167.0608 LAYER C4 ;
    ANTENNADIFFAREA 167.0608 LAYER C3 ;
    ANTENNADIFFAREA 167.0608 LAYER C5 ;
    ANTENNADIFFAREA 167.0608 LAYER JA ;
    ANTENNADIFFAREA 167.0608 LAYER QA ;
    ANTENNADIFFAREA 167.0608 LAYER QB ;
    ANTENNADIFFAREA 167.0608 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
        RECT 2 24 58 28.8 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
    END
  END PAD_B
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.84 79.86 30.98 80 ;
    END
  END VDDQ
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C1 ;
      ANTENNAMAXAREACAR 59.65625 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.2 79.86 14.34 80 ;
    END
  END D_LVDS_I[1]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C1 ;
      ANTENNAMAXAREACAR 60.30625 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.84 79.86 17.98 80 ;
    END
  END D_LVDS_I[0]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.637946 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.68 79.86 39.82 80 ;
    END
  END D_IOSG_I[9]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.518659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.16 79.86 39.3 80 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.594022 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.64 79.86 38.78 80 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.369792 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.12 79.86 38.26 80 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.446458 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.6 79.86 37.74 80 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.136806 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.08 79.86 37.22 80 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.214583 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.56 79.86 36.7 80 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.670735 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.04 79.86 36.18 80 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.747794 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.52 79.86 35.66 80 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C1 ;
      ANTENNAMAXAREACAR 2.443131 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.8 79.86 42.94 80 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C1 ;
      ANTENNAMAXAREACAR 2.582738 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.28 79.86 42.42 80 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C1 ;
      ANTENNAMAXAREACAR 2.733211 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.76 79.86 41.9 80 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.179861 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.24 79.86 41.38 80 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.253194 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.72 79.86 40.86 80 ;
    END
  END D_IOSG_I[11]
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.32 79.86 30.46 80 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_RTERMCAL_LLHVT28_V

MACRO RIIO_EG1D80V_RTERMCAL_LVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_LVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.564137 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.2 79.86 40.34 80 ;
    END
  END D_IOSG_I[10]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2212 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.36 79.86 5.5 80 ;
    END
  END RESULT_O[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.84 79.86 4.98 80 ;
    END
  END RESULT_O[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.336729 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.4 79.86 19.54 80 ;
    END
  END MODE_I[1]
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.869565 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.04 79.86 23.18 80 ;
    END
  END MODE_I[0]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.058036 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.92 79.86 7.06 80 ;
    END
  END D_LVDS_I[3]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.736607 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.56 79.86 10.7 80 ;
    END
  END D_LVDS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 68.1725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 493.9475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 364.8 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 235.02 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.5176 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JV ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JW ;
    ANTENNAPARTIALCUTAREA 7.031552 LAYER A2 ;
    ANTENNADIFFAREA 167.0608 LAYER C4 ;
    ANTENNADIFFAREA 167.0608 LAYER C3 ;
    ANTENNADIFFAREA 167.0608 LAYER C5 ;
    ANTENNADIFFAREA 167.0608 LAYER JA ;
    ANTENNADIFFAREA 167.0608 LAYER QA ;
    ANTENNADIFFAREA 167.0608 LAYER QB ;
    ANTENNADIFFAREA 167.0608 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
        RECT 2 24 58 28.8 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
    END
  END PAD_B
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.84 79.86 30.98 80 ;
    END
  END VDDQ
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.450893 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.2 79.86 14.34 80 ;
    END
  END D_LVDS_I[1]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.129464 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.84 79.86 17.98 80 ;
    END
  END D_LVDS_I[0]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.637946 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.68 79.86 39.82 80 ;
    END
  END D_IOSG_I[9]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.518659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.16 79.86 39.3 80 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.594022 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.64 79.86 38.78 80 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.369792 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.12 79.86 38.26 80 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.446458 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.6 79.86 37.74 80 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.136806 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.08 79.86 37.22 80 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.214583 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.56 79.86 36.7 80 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.670735 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.04 79.86 36.18 80 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.747794 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.52 79.86 35.66 80 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C1 ;
      ANTENNAMAXAREACAR 2.443131 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.8 79.86 42.94 80 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C1 ;
      ANTENNAMAXAREACAR 2.582738 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.28 79.86 42.42 80 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C1 ;
      ANTENNAMAXAREACAR 2.733211 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.76 79.86 41.9 80 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.179861 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.24 79.86 41.38 80 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.253194 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.72 79.86 40.86 80 ;
    END
  END D_IOSG_I[11]
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.32 79.86 30.46 80 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_RTERMCAL_LVT28_V

MACRO RIIO_EG1D80V_RTERMCAL_RVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.564137 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.2 79.86 40.34 80 ;
    END
  END D_IOSG_I[10]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2212 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.36 79.86 5.5 80 ;
    END
  END RESULT_O[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.84 79.86 4.98 80 ;
    END
  END RESULT_O[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.336729 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.4 79.86 19.54 80 ;
    END
  END MODE_I[1]
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.869565 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.04 79.86 23.18 80 ;
    END
  END MODE_I[0]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.058036 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.92 79.86 7.06 80 ;
    END
  END D_LVDS_I[3]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.736607 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.56 79.86 10.7 80 ;
    END
  END D_LVDS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 68.1725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 493.9475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 364.8 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 235.02 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.5176 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JV ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JW ;
    ANTENNAPARTIALCUTAREA 7.031552 LAYER A2 ;
    ANTENNADIFFAREA 167.0608 LAYER C4 ;
    ANTENNADIFFAREA 167.0608 LAYER C3 ;
    ANTENNADIFFAREA 167.0608 LAYER C5 ;
    ANTENNADIFFAREA 167.0608 LAYER JA ;
    ANTENNADIFFAREA 167.0608 LAYER QA ;
    ANTENNADIFFAREA 167.0608 LAYER QB ;
    ANTENNADIFFAREA 167.0608 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
        RECT 2 24 58 28.8 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
    END
  END PAD_B
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.84 79.86 30.98 80 ;
    END
  END VDDQ
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.450893 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.2 79.86 14.34 80 ;
    END
  END D_LVDS_I[1]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.129464 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.84 79.86 17.98 80 ;
    END
  END D_LVDS_I[0]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.637946 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.68 79.86 39.82 80 ;
    END
  END D_IOSG_I[9]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.518659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.16 79.86 39.3 80 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.594022 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.64 79.86 38.78 80 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.369792 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.12 79.86 38.26 80 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.446458 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.6 79.86 37.74 80 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.136806 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.08 79.86 37.22 80 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.214583 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.56 79.86 36.7 80 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.670735 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.04 79.86 36.18 80 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.747794 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.52 79.86 35.66 80 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C1 ;
      ANTENNAMAXAREACAR 2.443131 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.8 79.86 42.94 80 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C1 ;
      ANTENNAMAXAREACAR 2.582738 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.28 79.86 42.42 80 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C1 ;
      ANTENNAMAXAREACAR 2.733211 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.76 79.86 41.9 80 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.179861 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.24 79.86 41.38 80 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.253194 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.72 79.86 40.86 80 ;
    END
  END D_IOSG_I[11]
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.32 79.86 30.46 80 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_RTERMCAL_RVT28_V

MACRO RIIO_EG1D80V_RTERMCAL_SLVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_SLVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.564137 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.2 79.86 40.34 80 ;
    END
  END D_IOSG_I[10]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2212 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.36 79.86 5.5 80 ;
    END
  END RESULT_O[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.84 79.86 4.98 80 ;
    END
  END RESULT_O[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.336729 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.4 79.86 19.54 80 ;
    END
  END MODE_I[1]
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.869565 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.04 79.86 23.18 80 ;
    END
  END MODE_I[0]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.058036 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.92 79.86 7.06 80 ;
    END
  END D_LVDS_I[3]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.736607 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.56 79.86 10.7 80 ;
    END
  END D_LVDS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
    END
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 68.1725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 493.9475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 364.8 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 235.02 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.5176 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JV ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JW ;
    ANTENNAPARTIALCUTAREA 7.031552 LAYER A2 ;
    ANTENNADIFFAREA 167.0608 LAYER C4 ;
    ANTENNADIFFAREA 167.0608 LAYER C3 ;
    ANTENNADIFFAREA 167.0608 LAYER C5 ;
    ANTENNADIFFAREA 167.0608 LAYER JA ;
    ANTENNADIFFAREA 167.0608 LAYER QA ;
    ANTENNADIFFAREA 167.0608 LAYER QB ;
    ANTENNADIFFAREA 167.0608 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
        RECT 2 24 58 28.8 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
    END
  END PAD_B
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.84 79.86 30.98 80 ;
    END
  END VDDQ
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.450893 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.2 79.86 14.34 80 ;
    END
  END D_LVDS_I[1]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.129464 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.84 79.86 17.98 80 ;
    END
  END D_LVDS_I[0]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.637946 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.68 79.86 39.82 80 ;
    END
  END D_IOSG_I[9]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.518659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.16 79.86 39.3 80 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.594022 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.64 79.86 38.78 80 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.369792 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.12 79.86 38.26 80 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.446458 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.6 79.86 37.74 80 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.136806 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.08 79.86 37.22 80 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.214583 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.56 79.86 36.7 80 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.670735 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.04 79.86 36.18 80 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.747794 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.52 79.86 35.66 80 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C1 ;
      ANTENNAMAXAREACAR 2.443131 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.8 79.86 42.94 80 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C1 ;
      ANTENNAMAXAREACAR 2.582738 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.28 79.86 42.42 80 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C1 ;
      ANTENNAMAXAREACAR 2.733211 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.76 79.86 41.9 80 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.179861 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.24 79.86 41.38 80 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.253194 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.72 79.86 40.86 80 ;
    END
  END D_IOSG_I[11]
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.32 79.86 30.46 80 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_RTERMCAL_SLVT28_V


MACRO RIIO_EG1D80V_HPLVDS_RX_SLVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_HPLVDS_RX_SLVT28_H 0 0 ;
  SIZE 80 BY 180 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN A_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 585.0375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1004.7775 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1090.5675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 609.1608 LAYER JA ;
    ANTENNAPARTIALMETALAREA 1285.0008 LAYER QA ;
    ANTENNAPARTIALMETALAREA 615.8808 LAYER QB ;
    ANTENNAPARTIALMETALAREA 296.94 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 14.911072 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 17.86928 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 33.42222 LAYER YS ;
    ANTENNAPARTIALCUTAREA 69.12 LAYER JV ;
    ANTENNAPARTIALCUTAREA 69.12 LAYER JW ;
    ANTENNAPARTIALCUTAREA 10.117536 LAYER A2 ;
    ANTENNADIFFAREA 153.2196 LAYER C4 ;
    ANTENNADIFFAREA 153.2196 LAYER C3 ;
    ANTENNADIFFAREA 153.2196 LAYER C5 ;
    ANTENNADIFFAREA 153.2196 LAYER JA ;
    ANTENNADIFFAREA 153.2196 LAYER QA ;
    ANTENNADIFFAREA 153.2196 LAYER QB ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 87.6 ;
        RECT 0 0.8 2.4 5.6 ;
        RECT 0 7 2.4 11.8 ;
        RECT 0 13.2 2.4 18 ;
        RECT 0 19.4 2.4 24.2 ;
        RECT 0 25.6 2.4 30.4 ;
        RECT 0 31.8 2.4 36.6 ;
        RECT 0 38 2.4 42.8 ;
        RECT 0 44.2 2.4 49 ;
        RECT 0 50.4 2.4 55.2 ;
        RECT 0 56.6 2.4 61.4 ;
        RECT 0 62.8 2.4 67.6 ;
        RECT 0 69 2.4 73.8 ;
        RECT 0 75.2 2.4 80 ;
        RECT 0 81.4 2.4 86.2 ;
      LAYER QA ;
        RECT 0 0.8 2.4 5.6 ;
        RECT 0 7 2.4 11.8 ;
        RECT 0 13.2 2.4 18 ;
        RECT 0 19.4 2.4 24.2 ;
        RECT 0 25.6 2.4 30.4 ;
        RECT 0 31.8 2.4 36.6 ;
        RECT 0 38 2.4 42.8 ;
        RECT 0 44.2 2.4 49 ;
        RECT 0 50.4 2.4 55.2 ;
        RECT 0 56.6 2.4 61.4 ;
        RECT 0 62.8 2.4 67.6 ;
        RECT 0 69 2.4 73.8 ;
        RECT 0 75.2 2.4 80 ;
        RECT 0 81.4 2.4 86.2 ;
      LAYER C2 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER C3 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER C4 ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 99.95 1.85 103.55 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER JA ;
        RECT 0 0.8 2.4 5.6 ;
        RECT 0 7 2.4 11.8 ;
        RECT 0 13.2 2.4 18 ;
        RECT 0 19.4 2.4 24.2 ;
        RECT 0 25.6 2.4 30.4 ;
        RECT 0 31.8 2.4 36.6 ;
        RECT 0 38 2.4 42.8 ;
        RECT 0 44.2 2.4 49 ;
        RECT 0 50.4 2.4 55.2 ;
        RECT 0 56.6 2.4 61.4 ;
        RECT 0 62.8 2.4 67.6 ;
        RECT 0 69 2.4 73.8 ;
        RECT 0 75.2 2.4 80 ;
        RECT 0 81.4 2.4 86.2 ;
      LAYER C5 ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 99.95 1.85 103.55 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
    END
  END A_PAD_B
  PIN RX_GAIN_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8955 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 347.558333 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 86.67 80 86.83 ;
    END
  END RX_GAIN_I[1]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 180 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 180 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 168.2 80 173 ;
      LAYER QA ;
        RECT 75.2 168.2 80 173 ;
      LAYER JA ;
        RECT 75.2 168.2 80 173 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 155.8 80 160.6 ;
      LAYER QA ;
        RECT 75.2 155.8 80 160.6 ;
      LAYER JA ;
        RECT 75.2 155.8 80 160.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 143.4 80 148.2 ;
      LAYER QA ;
        RECT 75.2 143.4 80 148.2 ;
      LAYER JA ;
        RECT 75.2 143.4 80 148.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 131 80 135.8 ;
      LAYER QA ;
        RECT 75.2 131 80 135.8 ;
      LAYER JA ;
        RECT 75.2 131 80 135.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 118.6 80 123.4 ;
      LAYER QA ;
        RECT 75.2 118.6 80 123.4 ;
      LAYER JA ;
        RECT 75.2 118.6 80 123.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 106.2 80 111 ;
      LAYER QA ;
        RECT 75.2 106.2 80 111 ;
      LAYER JA ;
        RECT 75.2 106.2 80 111 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 93.8 80 98.6 ;
      LAYER QA ;
        RECT 75.2 93.8 80 98.6 ;
      LAYER JA ;
        RECT 75.2 93.8 80 98.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 81.4 80 86.2 ;
      LAYER QA ;
        RECT 75.2 81.4 80 86.2 ;
      LAYER JA ;
        RECT 75.2 81.4 80 86.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 69 80 73.8 ;
      LAYER QA ;
        RECT 75.2 69 80 73.8 ;
      LAYER JA ;
        RECT 75.2 69 80 73.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 56.6 80 61.4 ;
      LAYER QA ;
        RECT 75.2 56.6 80 61.4 ;
      LAYER JA ;
        RECT 75.2 56.6 80 61.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 44.2 80 49 ;
      LAYER QA ;
        RECT 75.2 44.2 80 49 ;
      LAYER JA ;
        RECT 75.2 44.2 80 49 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 31.8 80 36.6 ;
      LAYER QA ;
        RECT 75.2 31.8 80 36.6 ;
      LAYER JA ;
        RECT 75.2 31.8 80 36.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 19.4 80 24.2 ;
      LAYER QA ;
        RECT 75.2 19.4 80 24.2 ;
      LAYER JA ;
        RECT 75.2 19.4 80 24.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 7 80 11.8 ;
      LAYER QA ;
        RECT 75.2 7 80 11.8 ;
      LAYER JA ;
        RECT 75.2 7 80 11.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 180 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 180 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 180 ;
    END
  END VDDIO
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.408 LAYER C4 ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER C4 ;
        RECT 39.575 0 40.825 180 ;
    END
  END VBIAS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 180 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 180 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 180 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 180 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 180 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 174.4 80 179.2 ;
      LAYER QA ;
        RECT 75.2 174.4 80 179.2 ;
      LAYER JA ;
        RECT 75.2 174.4 80 179.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 162 80 166.8 ;
      LAYER QA ;
        RECT 75.2 162 80 166.8 ;
      LAYER JA ;
        RECT 75.2 162 80 166.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 149.6 80 154.4 ;
      LAYER QA ;
        RECT 75.2 149.6 80 154.4 ;
      LAYER JA ;
        RECT 75.2 149.6 80 154.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 137.2 80 142 ;
      LAYER QA ;
        RECT 75.2 137.2 80 142 ;
      LAYER JA ;
        RECT 75.2 137.2 80 142 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 124.8 80 129.6 ;
      LAYER QA ;
        RECT 75.2 124.8 80 129.6 ;
      LAYER JA ;
        RECT 75.2 124.8 80 129.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 112.4 80 117.2 ;
      LAYER QA ;
        RECT 75.2 112.4 80 117.2 ;
      LAYER JA ;
        RECT 75.2 112.4 80 117.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 100 80 104.8 ;
      LAYER QA ;
        RECT 75.2 100 80 104.8 ;
      LAYER JA ;
        RECT 75.2 100 80 104.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 87.6 80 92.4 ;
      LAYER QA ;
        RECT 75.2 87.6 80 92.4 ;
      LAYER JA ;
        RECT 75.2 87.6 80 92.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 75.2 80 80 ;
      LAYER QA ;
        RECT 75.2 75.2 80 80 ;
      LAYER JA ;
        RECT 75.2 75.2 80 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 62.8 80 67.6 ;
      LAYER QA ;
        RECT 75.2 62.8 80 67.6 ;
      LAYER JA ;
        RECT 75.2 62.8 80 67.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 50.4 80 55.2 ;
      LAYER QA ;
        RECT 75.2 50.4 80 55.2 ;
      LAYER JA ;
        RECT 75.2 50.4 80 55.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 38 80 42.8 ;
      LAYER QA ;
        RECT 75.2 38 80 42.8 ;
      LAYER JA ;
        RECT 75.2 38 80 42.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 25.6 80 30.4 ;
      LAYER QA ;
        RECT 75.2 25.6 80 30.4 ;
      LAYER JA ;
        RECT 75.2 25.6 80 30.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 13.2 80 18 ;
      LAYER QA ;
        RECT 75.2 13.2 80 18 ;
      LAYER JA ;
        RECT 75.2 13.2 80 18 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 0.8 80 5.6 ;
      LAYER QA ;
        RECT 75.2 0.8 80 5.6 ;
      LAYER JA ;
        RECT 75.2 0.8 80 5.6 ;
    END
  END VSS
  PIN RX_CTLE_RES_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7195 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.639394 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 91.09 80 91.25 ;
    END
  END RX_CTLE_RES_I[2]
  PIN EI_DETECT_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2128 LAYER C2 ;
    ANTENNADIFFAREA 0.081 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 49.23 80 49.39 ;
    END
  END EI_DETECT_O
  PIN EI_DETECT_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 35.102484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 131.91 80 132.07 ;
    END
  END EI_DETECT_EN_I
  PIN RTERM_TRIM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 177.15 80 177.31 ;
    END
  END RTERM_TRIM_I[3]
  PIN B_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1022.5375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1004.7775 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1090.5675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 609.12 LAYER JA ;
    ANTENNAPARTIALMETALAREA 1284.96 LAYER QA ;
    ANTENNAPARTIALMETALAREA 615.84 LAYER QB ;
    ANTENNAPARTIALMETALAREA 747.92 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 19.085088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 17.86928 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 33.42222 LAYER YS ;
    ANTENNAPARTIALCUTAREA 69.12 LAYER JV ;
    ANTENNAPARTIALCUTAREA 69.12 LAYER JW ;
    ANTENNAPARTIALCUTAREA 10.713824 LAYER A2 ;
    ANTENNADIFFAREA 153.2196 LAYER C4 ;
    ANTENNADIFFAREA 153.2196 LAYER C3 ;
    ANTENNADIFFAREA 153.2196 LAYER C5 ;
    ANTENNADIFFAREA 153.2196 LAYER JA ;
    ANTENNADIFFAREA 153.2196 LAYER QA ;
    ANTENNADIFFAREA 153.2196 LAYER QB ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 92.4 28.8 178 ;
        RECT 0 93.817 2.4 98.617 ;
        RECT 0 100.017 2.4 104.817 ;
        RECT 0 106.217 2.4 111.017 ;
        RECT 0 112.417 2.4 117.217 ;
        RECT 0 118.617 2.4 123.417 ;
        RECT 0 124.817 2.4 129.617 ;
        RECT 0 131.017 2.4 135.817 ;
        RECT 0 137.217 2.4 142.017 ;
        RECT 0 143.417 2.4 148.217 ;
        RECT 0 149.617 2.4 154.417 ;
        RECT 0 155.817 2.4 160.617 ;
        RECT 0 162.017 2.4 166.817 ;
        RECT 0 168.217 2.4 173.017 ;
        RECT 0 174.417 2.4 179.217 ;
      LAYER QA ;
        RECT 0 93.817 2.4 98.617 ;
        RECT 0 100.017 2.4 104.817 ;
        RECT 0 106.217 2.4 111.017 ;
        RECT 0 112.417 2.4 117.217 ;
        RECT 0 118.617 2.4 123.417 ;
        RECT 0 124.817 2.4 129.617 ;
        RECT 0 131.017 2.4 135.817 ;
        RECT 0 137.217 2.4 142.017 ;
        RECT 0 143.417 2.4 148.217 ;
        RECT 0 149.617 2.4 154.417 ;
        RECT 0 155.817 2.4 160.617 ;
        RECT 0 162.017 2.4 166.817 ;
        RECT 0 168.217 2.4 173.017 ;
        RECT 0 174.417 2.4 179.217 ;
      LAYER C2 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
      LAYER C3 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
      LAYER C4 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
        RECT 0 76.45 1.85 80.05 ;
        RECT 0 81.15 1.85 84.75 ;
      LAYER JA ;
        RECT 0 93.817 2.4 98.617 ;
        RECT 0 100.017 2.4 104.817 ;
        RECT 0 106.217 2.4 111.017 ;
        RECT 0 112.417 2.4 117.217 ;
        RECT 0 118.617 2.4 123.417 ;
        RECT 0 124.817 2.4 129.617 ;
        RECT 0 131.017 2.4 135.817 ;
        RECT 0 137.217 2.4 142.017 ;
        RECT 0 143.417 2.4 148.217 ;
        RECT 0 149.617 2.4 154.417 ;
        RECT 0 155.817 2.4 160.617 ;
        RECT 0 162.017 2.4 166.817 ;
        RECT 0 168.217 2.4 173.017 ;
        RECT 0 174.417 2.4 179.217 ;
      LAYER C5 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
        RECT 0 76.45 1.85 80.05 ;
        RECT 0 81.15 1.85 84.75 ;
    END
  END B_PAD_B
  PIN RTERM_TRIM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 176.63 80 176.79 ;
    END
  END RTERM_TRIM_I[2]
  PIN RTERM_TRIM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 176.11 80 176.27 ;
    END
  END RTERM_TRIM_I[1]
  PIN RTERM_TRIM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 175.59 80 175.75 ;
    END
  END RTERM_TRIM_I[0]
  PIN RTERM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 28.891274 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 175.07 80 175.23 ;
    END
  END RTERM_EN_I
  PIN RX_CTLE_CAP_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7195 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 463.455556 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 88.75 80 88.91 ;
    END
  END RX_CTLE_CAP_I[2]
  PIN RX_GAIN_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8515 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 347.915 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 87.19 80 87.35 ;
    END
  END RX_GAIN_I[2]
  PIN DI_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2128 LAYER C2 ;
    ANTENNADIFFAREA 0.16192 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 129.83 80 129.99 ;
    END
  END DI_O
  PIN RX_CTLE_RES_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8515 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.287879 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 92.65 80 92.81 ;
    END
  END RX_CTLE_RES_I[5]
  PIN RX_CTLE_RES_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8955 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 471.867677 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 93.17 80 93.33 ;
    END
  END RX_CTLE_RES_I[6]
  PIN RX_GAIN_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8075 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 346.412778 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 87.71 80 87.87 ;
    END
  END RX_GAIN_I[3]
  PIN RX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C2 ;
      ANTENNAMAXAREACAR 56.869643 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 128.27 80 128.43 ;
    END
  END RX_POL_I
  PIN RX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 35.102484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 132.95 80 133.11 ;
    END
  END RX_VCM_EN_I
  PIN RX_CTLE_RES_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7635 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.522222 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 91.61 80 91.77 ;
    END
  END RX_CTLE_RES_I[3]
  PIN RX_CTLE_RES_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8075 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.405051 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 92.13 80 92.29 ;
    END
  END RX_CTLE_RES_I[4]
  PIN RX_CTLE_RES_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9395 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 473.457576 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 93.69 80 93.85 ;
    END
  END RX_CTLE_RES_I[7]
  PIN RX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9395 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 346.633889 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 86.15 80 86.31 ;
    END
  END RX_EN_I
  PIN RX_CTLE_CAP_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6755 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 478.89798 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 89.27 80 89.43 ;
    END
  END RX_CTLE_CAP_I[3]
  PIN RX_CTLE_RES_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6755 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.756566 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 90.57 80 90.73 ;
    END
  END RX_CTLE_RES_I[1]
  PIN RX_CTLE_CAP_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7635 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 468.536364 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 88.23 80 88.39 ;
    END
  END RX_CTLE_CAP_I[1]
  OBS
    LAYER CA ;
      RECT 0 0 80 180 ;
    LAYER M1 ;
      RECT 0 0 80 180 ;
    LAYER V1 ;
      RECT 0 0 80 180 ;
    LAYER M2 ;
      RECT 0 0 80 180 ;
    LAYER A1 ;
      RECT 0 0 80 180 ;
    LAYER C2 ;
      RECT 0 0 80 180 ;
    LAYER CB ;
      RECT 0 0 80 180 ;
    LAYER JV ;
      RECT 0 0 80 180 ;
    LAYER YS ;
      RECT 0 0 80 180 ;
    LAYER JW ;
      RECT 0 0 80 180 ;
    LAYER QB ;
      RECT 0 0 80 180 ;
    LAYER QA ;
      RECT 0 0 80 180 ;
    LAYER JA ;
      RECT 0 0 80 180 ;
    LAYER AY ;
      RECT 0 0 80 180 ;
    LAYER C1 ;
      RECT 0 0 80 180 ;
    LAYER C5 ;
      RECT 0 0 80 180 ;
    LAYER C4 ;
      RECT 0 0 80 180 ;
    LAYER C3 ;
      RECT 0 0 80 180 ;
    LAYER A4 ;
      RECT 0 0 80 180 ;
    LAYER A3 ;
      RECT 0 0 80 180 ;
    LAYER A2 ;
      RECT 0 0 80 180 ;
  END
END RIIO_EG1D80V_HPLVDS_RX_SLVT28_H

MACRO RIIO_EG1D80V_HPLVDS_TX_SLVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_HPLVDS_TX_SLVT28_H 0 0 ;
  SIZE 80 BY 180 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN A_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 585.0375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1004.7775 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1090.5675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 609.1608 LAYER JA ;
    ANTENNAPARTIALMETALAREA 1285.0008 LAYER QA ;
    ANTENNAPARTIALMETALAREA 615.8808 LAYER QB ;
    ANTENNAPARTIALMETALAREA 296.94 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 14.911072 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 17.86928 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 33.42222 LAYER YS ;
    ANTENNAPARTIALCUTAREA 69.12 LAYER JV ;
    ANTENNAPARTIALCUTAREA 69.12 LAYER JW ;
    ANTENNAPARTIALCUTAREA 10.117536 LAYER A2 ;
    ANTENNADIFFAREA 206.9796 LAYER C4 ;
    ANTENNADIFFAREA 206.9796 LAYER C3 ;
    ANTENNADIFFAREA 206.9796 LAYER C5 ;
    ANTENNADIFFAREA 206.9796 LAYER JA ;
    ANTENNADIFFAREA 206.9796 LAYER QA ;
    ANTENNADIFFAREA 206.9796 LAYER QB ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 87.6 ;
        RECT 0 0.8 2.4 5.6 ;
        RECT 0 7 2.4 11.8 ;
        RECT 0 13.2 2.4 18 ;
        RECT 0 19.4 2.4 24.2 ;
        RECT 0 25.6 2.4 30.4 ;
        RECT 0 31.8 2.4 36.6 ;
        RECT 0 38 2.4 42.8 ;
        RECT 0 44.2 2.4 49 ;
        RECT 0 50.4 2.4 55.2 ;
        RECT 0 56.6 2.4 61.4 ;
        RECT 0 62.8 2.4 67.6 ;
        RECT 0 69 2.4 73.8 ;
        RECT 0 75.2 2.4 80 ;
        RECT 0 81.4 2.4 86.2 ;
      LAYER QA ;
        RECT 0 0.8 2.4 5.6 ;
        RECT 0 7 2.4 11.8 ;
        RECT 0 13.2 2.4 18 ;
        RECT 0 19.4 2.4 24.2 ;
        RECT 0 25.6 2.4 30.4 ;
        RECT 0 31.8 2.4 36.6 ;
        RECT 0 38 2.4 42.8 ;
        RECT 0 44.2 2.4 49 ;
        RECT 0 50.4 2.4 55.2 ;
        RECT 0 56.6 2.4 61.4 ;
        RECT 0 62.8 2.4 67.6 ;
        RECT 0 69 2.4 73.8 ;
        RECT 0 75.2 2.4 80 ;
        RECT 0 81.4 2.4 86.2 ;
      LAYER C2 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER C3 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER C4 ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 99.95 1.85 103.55 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER JA ;
        RECT 0 0.8 2.4 5.6 ;
        RECT 0 7 2.4 11.8 ;
        RECT 0 13.2 2.4 18 ;
        RECT 0 19.4 2.4 24.2 ;
        RECT 0 25.6 2.4 30.4 ;
        RECT 0 31.8 2.4 36.6 ;
        RECT 0 38 2.4 42.8 ;
        RECT 0 44.2 2.4 49 ;
        RECT 0 50.4 2.4 55.2 ;
        RECT 0 56.6 2.4 61.4 ;
        RECT 0 62.8 2.4 67.6 ;
        RECT 0 69 2.4 73.8 ;
        RECT 0 75.2 2.4 80 ;
        RECT 0 81.4 2.4 86.2 ;
      LAYER C5 ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 99.95 1.85 103.55 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
    END
  END A_PAD_B
  PIN TX_FFE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23216 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02128 LAYER C2 ;
      ANTENNAMAXAREACAR 26.403195 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 129.31 80 129.47 ;
    END
  END TX_FFE_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 180 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 180 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 180 ;
    END
  END VDDIO
  PIN RX_GAIN_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8955 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 347.558333 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 86.67 80 86.83 ;
    END
  END RX_GAIN_I[1]
  PIN TX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C2 ;
      ANTENNAMAXAREACAR 54.698214 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 127.75 80 127.91 ;
    END
  END TX_POL_I
  PIN TX_EI_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0112 LAYER C2 ;
      ANTENNAMAXAREACAR 99.871429 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 128.79 80 128.95 ;
    END
  END TX_EI_I
  PIN TX_BIAS_OD_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 35.102484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 132.43 80 132.59 ;
    END
  END TX_BIAS_OD_I
  PIN TX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 28.164002 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 151.15 80 151.31 ;
    END
  END TX_EN_I
  PIN TX_BIAS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 153.23 80 153.39 ;
    END
  END TX_BIAS_I[3]
  PIN TX_VCM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 150.11 80 150.27 ;
    END
  END TX_VCM_I[2]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 180 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 180 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 180 ;
    END
  END VSSIO
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.408 LAYER C4 ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER C4 ;
        RECT 39.575 0 40.825 180 ;
    END
  END VBIAS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 180 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 180 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 168.2 80 173 ;
      LAYER QA ;
        RECT 75.2 168.2 80 173 ;
      LAYER JA ;
        RECT 75.2 168.2 80 173 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 155.8 80 160.6 ;
      LAYER QA ;
        RECT 75.2 155.8 80 160.6 ;
      LAYER JA ;
        RECT 75.2 155.8 80 160.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 143.4 80 148.2 ;
      LAYER QA ;
        RECT 75.2 143.4 80 148.2 ;
      LAYER JA ;
        RECT 75.2 143.4 80 148.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 131 80 135.8 ;
      LAYER QA ;
        RECT 75.2 131 80 135.8 ;
      LAYER JA ;
        RECT 75.2 131 80 135.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 118.6 80 123.4 ;
      LAYER QA ;
        RECT 75.2 118.6 80 123.4 ;
      LAYER JA ;
        RECT 75.2 118.6 80 123.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 106.2 80 111 ;
      LAYER QA ;
        RECT 75.2 106.2 80 111 ;
      LAYER JA ;
        RECT 75.2 106.2 80 111 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 93.8 80 98.6 ;
      LAYER QA ;
        RECT 75.2 93.8 80 98.6 ;
      LAYER JA ;
        RECT 75.2 93.8 80 98.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 81.4 80 86.2 ;
      LAYER QA ;
        RECT 75.2 81.4 80 86.2 ;
      LAYER JA ;
        RECT 75.2 81.4 80 86.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 69 80 73.8 ;
      LAYER QA ;
        RECT 75.2 69 80 73.8 ;
      LAYER JA ;
        RECT 75.2 69 80 73.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 56.6 80 61.4 ;
      LAYER QA ;
        RECT 75.2 56.6 80 61.4 ;
      LAYER JA ;
        RECT 75.2 56.6 80 61.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 44.2 80 49 ;
      LAYER QA ;
        RECT 75.2 44.2 80 49 ;
      LAYER JA ;
        RECT 75.2 44.2 80 49 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 31.8 80 36.6 ;
      LAYER QA ;
        RECT 75.2 31.8 80 36.6 ;
      LAYER JA ;
        RECT 75.2 31.8 80 36.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 19.4 80 24.2 ;
      LAYER QA ;
        RECT 75.2 19.4 80 24.2 ;
      LAYER JA ;
        RECT 75.2 19.4 80 24.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 7 80 11.8 ;
      LAYER QA ;
        RECT 75.2 7 80 11.8 ;
      LAYER JA ;
        RECT 75.2 7 80 11.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 180 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 180 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 174.4 80 179.2 ;
      LAYER QA ;
        RECT 75.2 174.4 80 179.2 ;
      LAYER JA ;
        RECT 75.2 174.4 80 179.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 162 80 166.8 ;
      LAYER QA ;
        RECT 75.2 162 80 166.8 ;
      LAYER JA ;
        RECT 75.2 162 80 166.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 149.6 80 154.4 ;
      LAYER QA ;
        RECT 75.2 149.6 80 154.4 ;
      LAYER JA ;
        RECT 75.2 149.6 80 154.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 137.2 80 142 ;
      LAYER QA ;
        RECT 75.2 137.2 80 142 ;
      LAYER JA ;
        RECT 75.2 137.2 80 142 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 124.8 80 129.6 ;
      LAYER QA ;
        RECT 75.2 124.8 80 129.6 ;
      LAYER JA ;
        RECT 75.2 124.8 80 129.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 112.4 80 117.2 ;
      LAYER QA ;
        RECT 75.2 112.4 80 117.2 ;
      LAYER JA ;
        RECT 75.2 112.4 80 117.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 100 80 104.8 ;
      LAYER QA ;
        RECT 75.2 100 80 104.8 ;
      LAYER JA ;
        RECT 75.2 100 80 104.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 87.6 80 92.4 ;
      LAYER QA ;
        RECT 75.2 87.6 80 92.4 ;
      LAYER JA ;
        RECT 75.2 87.6 80 92.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 75.2 80 80 ;
      LAYER QA ;
        RECT 75.2 75.2 80 80 ;
      LAYER JA ;
        RECT 75.2 75.2 80 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 62.8 80 67.6 ;
      LAYER QA ;
        RECT 75.2 62.8 80 67.6 ;
      LAYER JA ;
        RECT 75.2 62.8 80 67.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 50.4 80 55.2 ;
      LAYER QA ;
        RECT 75.2 50.4 80 55.2 ;
      LAYER JA ;
        RECT 75.2 50.4 80 55.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 38 80 42.8 ;
      LAYER QA ;
        RECT 75.2 38 80 42.8 ;
      LAYER JA ;
        RECT 75.2 38 80 42.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 25.6 80 30.4 ;
      LAYER QA ;
        RECT 75.2 25.6 80 30.4 ;
      LAYER JA ;
        RECT 75.2 25.6 80 30.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 13.2 80 18 ;
      LAYER QA ;
        RECT 75.2 13.2 80 18 ;
      LAYER JA ;
        RECT 75.2 13.2 80 18 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 0.8 80 5.6 ;
      LAYER QA ;
        RECT 75.2 0.8 80 5.6 ;
      LAYER JA ;
        RECT 75.2 0.8 80 5.6 ;
    END
  END VSS
  PIN RX_CTLE_RES_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7195 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.639394 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 91.09 80 91.25 ;
    END
  END RX_CTLE_RES_I[2]
  PIN TX_VCM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 149.59 80 149.75 ;
    END
  END TX_VCM_I[1]
  PIN EI_DETECT_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2128 LAYER C2 ;
    ANTENNADIFFAREA 0.081 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 49.23 80 49.39 ;
    END
  END EI_DETECT_O
  PIN EI_DETECT_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 35.102484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 131.91 80 132.07 ;
    END
  END EI_DETECT_EN_I
  PIN RTERM_TRIM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 177.15 80 177.31 ;
    END
  END RTERM_TRIM_I[3]
  PIN B_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1022.5375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1004.7775 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1090.5675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 609.12 LAYER JA ;
    ANTENNAPARTIALMETALAREA 1284.96 LAYER QA ;
    ANTENNAPARTIALMETALAREA 615.84 LAYER QB ;
    ANTENNAPARTIALMETALAREA 747.92 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 19.085088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 17.86928 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 33.42222 LAYER YS ;
    ANTENNAPARTIALCUTAREA 69.12 LAYER JV ;
    ANTENNAPARTIALCUTAREA 69.12 LAYER JW ;
    ANTENNAPARTIALCUTAREA 10.713824 LAYER A2 ;
    ANTENNADIFFAREA 206.9796 LAYER C4 ;
    ANTENNADIFFAREA 206.9796 LAYER C3 ;
    ANTENNADIFFAREA 206.9796 LAYER C5 ;
    ANTENNADIFFAREA 206.9796 LAYER JA ;
    ANTENNADIFFAREA 206.9796 LAYER QA ;
    ANTENNADIFFAREA 206.9796 LAYER QB ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 92.4 28.8 178 ;
        RECT 0 93.817 2.4 98.617 ;
        RECT 0 100.017 2.4 104.817 ;
        RECT 0 106.217 2.4 111.017 ;
        RECT 0 112.417 2.4 117.217 ;
        RECT 0 118.617 2.4 123.417 ;
        RECT 0 124.817 2.4 129.617 ;
        RECT 0 131.017 2.4 135.817 ;
        RECT 0 137.217 2.4 142.017 ;
        RECT 0 143.417 2.4 148.217 ;
        RECT 0 149.617 2.4 154.417 ;
        RECT 0 155.817 2.4 160.617 ;
        RECT 0 162.017 2.4 166.817 ;
        RECT 0 168.217 2.4 173.017 ;
        RECT 0 174.417 2.4 179.217 ;
      LAYER QA ;
        RECT 0 93.817 2.4 98.617 ;
        RECT 0 100.017 2.4 104.817 ;
        RECT 0 106.217 2.4 111.017 ;
        RECT 0 112.417 2.4 117.217 ;
        RECT 0 118.617 2.4 123.417 ;
        RECT 0 124.817 2.4 129.617 ;
        RECT 0 131.017 2.4 135.817 ;
        RECT 0 137.217 2.4 142.017 ;
        RECT 0 143.417 2.4 148.217 ;
        RECT 0 149.617 2.4 154.417 ;
        RECT 0 155.817 2.4 160.617 ;
        RECT 0 162.017 2.4 166.817 ;
        RECT 0 168.217 2.4 173.017 ;
        RECT 0 174.417 2.4 179.217 ;
      LAYER C2 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
      LAYER C3 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
      LAYER C4 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
        RECT 0 76.45 1.85 80.05 ;
        RECT 0 81.15 1.85 84.75 ;
      LAYER JA ;
        RECT 0 93.817 2.4 98.617 ;
        RECT 0 100.017 2.4 104.817 ;
        RECT 0 106.217 2.4 111.017 ;
        RECT 0 112.417 2.4 117.217 ;
        RECT 0 118.617 2.4 123.417 ;
        RECT 0 124.817 2.4 129.617 ;
        RECT 0 131.017 2.4 135.817 ;
        RECT 0 137.217 2.4 142.017 ;
        RECT 0 143.417 2.4 148.217 ;
        RECT 0 149.617 2.4 154.417 ;
        RECT 0 155.817 2.4 160.617 ;
        RECT 0 162.017 2.4 166.817 ;
        RECT 0 168.217 2.4 173.017 ;
        RECT 0 174.417 2.4 179.217 ;
      LAYER C5 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
        RECT 0 76.45 1.85 80.05 ;
        RECT 0 81.15 1.85 84.75 ;
    END
  END B_PAD_B
  PIN RTERM_TRIM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 176.63 80 176.79 ;
    END
  END RTERM_TRIM_I[2]
  PIN RTERM_TRIM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 176.11 80 176.27 ;
    END
  END RTERM_TRIM_I[1]
  PIN RTERM_TRIM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 175.59 80 175.75 ;
    END
  END RTERM_TRIM_I[0]
  PIN RTERM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 28.891274 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 175.07 80 175.23 ;
    END
  END RTERM_EN_I
  PIN RX_CTLE_CAP_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7195 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 463.455556 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 88.75 80 88.91 ;
    END
  END RX_CTLE_CAP_I[2]
  PIN RX_GAIN_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8515 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 347.915 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 87.19 80 87.35 ;
    END
  END RX_GAIN_I[2]
  PIN TX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 32.20556 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 148.55 80 148.71 ;
    END
  END TX_VCM_EN_I
  PIN TX_VCM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 150.63 80 150.79 ;
    END
  END TX_VCM_I[3]
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2128 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C2 ;
      ANTENNAMAXAREACAR 30.536607 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 130.87 80 131.03 ;
    END
  END DO_I
  PIN DI_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2128 LAYER C2 ;
    ANTENNADIFFAREA 0.16192 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 129.83 80 129.99 ;
    END
  END DI_O
  PIN RX_CTLE_RES_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8515 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.287879 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 92.65 80 92.81 ;
    END
  END RX_CTLE_RES_I[5]
  PIN RX_CTLE_RES_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8955 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 471.867677 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 93.17 80 93.33 ;
    END
  END RX_CTLE_RES_I[6]
  PIN TX_BIAS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 152.71 80 152.87 ;
    END
  END TX_BIAS_I[2]
  PIN RX_GAIN_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8075 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 346.412778 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 87.71 80 87.87 ;
    END
  END RX_GAIN_I[3]
  PIN RX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C2 ;
      ANTENNAMAXAREACAR 56.869643 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 128.27 80 128.43 ;
    END
  END RX_POL_I
  PIN RX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 35.102484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 132.95 80 133.11 ;
    END
  END RX_VCM_EN_I
  PIN TX_BIAS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 152.19 80 152.35 ;
    END
  END TX_BIAS_I[1]
  PIN RX_CTLE_RES_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7635 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.522222 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 91.61 80 91.77 ;
    END
  END RX_CTLE_RES_I[3]
  PIN RX_CTLE_RES_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8075 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.405051 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 92.13 80 92.29 ;
    END
  END RX_CTLE_RES_I[4]
  PIN TX_VCM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 149.07 80 149.23 ;
    END
  END TX_VCM_I[0]
  PIN TX_BIAS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 151.67 80 151.83 ;
    END
  END TX_BIAS_I[0]
  PIN RX_CTLE_RES_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9395 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 473.457576 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 93.69 80 93.85 ;
    END
  END RX_CTLE_RES_I[7]
  PIN RX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9395 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 346.633889 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 86.15 80 86.31 ;
    END
  END RX_EN_I
  PIN RX_CTLE_CAP_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6755 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 478.89798 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 89.27 80 89.43 ;
    END
  END RX_CTLE_CAP_I[3]
  PIN RX_CTLE_RES_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6755 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.756566 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 90.57 80 90.73 ;
    END
  END RX_CTLE_RES_I[1]
  PIN RX_CTLE_CAP_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7635 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 468.536364 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 88.23 80 88.39 ;
    END
  END RX_CTLE_CAP_I[1]
  OBS
    LAYER CA ;
      RECT 0 0 80 180 ;
    LAYER M1 ;
      RECT 0 0 80 180 ;
    LAYER V1 ;
      RECT 0 0 80 180 ;
    LAYER M2 ;
      RECT 0 0 80 180 ;
    LAYER A1 ;
      RECT 0 0 80 180 ;
    LAYER C2 ;
      RECT 0 0 80 180 ;
    LAYER CB ;
      RECT 0 0 80 180 ;
    LAYER JV ;
      RECT 0 0 80 180 ;
    LAYER YS ;
      RECT 0 0 80 180 ;
    LAYER JW ;
      RECT 0 0 80 180 ;
    LAYER QB ;
      RECT 0 0 80 180 ;
    LAYER QA ;
      RECT 0 0 80 180 ;
    LAYER JA ;
      RECT 0 0 80 180 ;
    LAYER AY ;
      RECT 0 0 80 180 ;
    LAYER C1 ;
      RECT 0 0 80 180 ;
    LAYER C5 ;
      RECT 0 0 80 180 ;
    LAYER C4 ;
      RECT 0 0 80 180 ;
    LAYER C3 ;
      RECT 0 0 80 180 ;
    LAYER A4 ;
      RECT 0 0 80 180 ;
    LAYER A3 ;
      RECT 0 0 80 180 ;
    LAYER A2 ;
      RECT 0 0 80 180 ;
  END
END RIIO_EG1D80V_HPLVDS_TX_SLVT28_H

MACRO RIIO_EG1D80V_RTERMCAL_HVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_HVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.46 80 40.6 ;
    END
  END VSSQ
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 567.2075 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 487.68 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 310.30352 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JV ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JW ;
    ANTENNAPARTIALCUTAREA 17.131488 LAYER A2 ;
    ANTENNADIFFAREA 152.2484 LAYER C4 ;
    ANTENNADIFFAREA 152.2484 LAYER C3 ;
    ANTENNADIFFAREA 152.2484 LAYER C5 ;
    ANTENNADIFFAREA 152.2484 LAYER JA ;
    ANTENNADIFFAREA 152.2484 LAYER QA ;
    ANTENNADIFFAREA 152.2484 LAYER QB ;
    ANTENNADIFFAREA 152.2484 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 98.217391 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.74 80 47.88 ;
    END
  END MODE_I[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 52.609456 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.22 80 47.36 ;
    END
  END MODE_I[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.7 80 46.84 ;
    END
  END RESULT_O[0]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.18 80 46.32 ;
    END
  END RESULT_O[1]
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.02 80 55.16 ;
    END
  END D_IOSG_I[10]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.811972 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.54 80 55.68 ;
    END
  END D_IOSG_I[11]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.82975 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.06 80 56.2 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C2 ;
      ANTENNAMAXAREACAR 14.865466 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.58 80 56.72 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C2 ;
      ANTENNAMAXAREACAR 14.455976 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.1 80 57.24 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C2 ;
      ANTENNAMAXAREACAR 13.688986 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.62 80 57.76 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.665245 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.34 80 50.48 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.666814 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.86 80 51 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.38 80 51.52 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.9 80 52.04 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.42 80 52.56 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.94 80 53.08 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.46 80 53.6 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.98 80 54.12 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 54.5 80 54.64 ;
    END
  END D_IOSG_I[9]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.629464 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.82 80 49.96 ;
    END
  END D_LVDS_I[0]
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.950893 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.3 80 49.44 ;
    END
  END D_LVDS_I[1]
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.98 80 41.12 ;
    END
  END VDDQ
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.236607 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.78 80 48.92 ;
    END
  END D_LVDS_I[2]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.558036 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.26 80 48.4 ;
    END
  END D_LVDS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_RTERMCAL_HVT28_H

MACRO RIIO_EG1D80V_RTERMCAL_LLHVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_LLHVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.46 80 40.6 ;
    END
  END VSSQ
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 567.2075 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 487.68 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 310.30352 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JV ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JW ;
    ANTENNAPARTIALCUTAREA 17.131488 LAYER A2 ;
    ANTENNADIFFAREA 152.2484 LAYER C4 ;
    ANTENNADIFFAREA 152.2484 LAYER C3 ;
    ANTENNADIFFAREA 152.2484 LAYER C5 ;
    ANTENNADIFFAREA 152.2484 LAYER JA ;
    ANTENNADIFFAREA 152.2484 LAYER QA ;
    ANTENNADIFFAREA 152.2484 LAYER QB ;
    ANTENNADIFFAREA 152.2484 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0184 LAYER C2 ;
      ANTENNAMAXAREACAR 138.063043 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.74 80 47.88 ;
    END
  END MODE_I[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.044 LAYER C2 ;
      ANTENNAMAXAREACAR 72.110568 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.22 80 47.36 ;
    END
  END MODE_I[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.03864 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.7 80 46.84 ;
    END
  END RESULT_O[0]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.03864 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.18 80 46.32 ;
    END
  END RESULT_O[1]
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.02 80 55.16 ;
    END
  END D_IOSG_I[10]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.811972 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.54 80 55.68 ;
    END
  END D_IOSG_I[11]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.82975 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.06 80 56.2 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C2 ;
      ANTENNAMAXAREACAR 14.865466 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.58 80 56.72 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C2 ;
      ANTENNAMAXAREACAR 14.455976 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.1 80 57.24 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C2 ;
      ANTENNAMAXAREACAR 13.688986 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.62 80 57.76 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.665245 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.34 80 50.48 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.666814 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.86 80 51 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.38 80 51.52 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.9 80 52.04 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.42 80 52.56 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.94 80 53.08 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.46 80 53.6 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.98 80 54.12 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 54.5 80 54.64 ;
    END
  END D_IOSG_I[9]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C2 ;
      ANTENNAMAXAREACAR 399.80625 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.82 80 49.96 ;
    END
  END D_LVDS_I[0]
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C2 ;
      ANTENNAMAXAREACAR 399.15625 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.3 80 49.44 ;
    END
  END D_LVDS_I[1]
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.98 80 41.12 ;
    END
  END VDDQ
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C2 ;
      ANTENNAMAXAREACAR 399.15625 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.78 80 48.92 ;
    END
  END D_LVDS_I[2]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C2 ;
      ANTENNAMAXAREACAR 399.15625 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.26 80 48.4 ;
    END
  END D_LVDS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_RTERMCAL_LLHVT28_H

MACRO RIIO_EG1D80V_RTERMCAL_LVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_LVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.46 80 40.6 ;
    END
  END VSSQ
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 567.2075 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 487.68 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 310.30352 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JV ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JW ;
    ANTENNAPARTIALCUTAREA 17.131488 LAYER A2 ;
    ANTENNADIFFAREA 152.2484 LAYER C4 ;
    ANTENNADIFFAREA 152.2484 LAYER C3 ;
    ANTENNADIFFAREA 152.2484 LAYER C5 ;
    ANTENNADIFFAREA 152.2484 LAYER JA ;
    ANTENNADIFFAREA 152.2484 LAYER QA ;
    ANTENNADIFFAREA 152.2484 LAYER QB ;
    ANTENNADIFFAREA 152.2484 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 98.217391 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.74 80 47.88 ;
    END
  END MODE_I[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 52.609456 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.22 80 47.36 ;
    END
  END MODE_I[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.7 80 46.84 ;
    END
  END RESULT_O[0]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.18 80 46.32 ;
    END
  END RESULT_O[1]
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.02 80 55.16 ;
    END
  END D_IOSG_I[10]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.811972 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.54 80 55.68 ;
    END
  END D_IOSG_I[11]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.82975 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.06 80 56.2 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C2 ;
      ANTENNAMAXAREACAR 14.865466 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.58 80 56.72 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C2 ;
      ANTENNAMAXAREACAR 14.455976 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.1 80 57.24 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C2 ;
      ANTENNAMAXAREACAR 13.688986 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.62 80 57.76 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.665245 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.34 80 50.48 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.666814 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.86 80 51 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.38 80 51.52 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.9 80 52.04 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.42 80 52.56 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.94 80 53.08 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.46 80 53.6 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.98 80 54.12 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 54.5 80 54.64 ;
    END
  END D_IOSG_I[9]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.629464 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.82 80 49.96 ;
    END
  END D_LVDS_I[0]
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.950893 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.3 80 49.44 ;
    END
  END D_LVDS_I[1]
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.98 80 41.12 ;
    END
  END VDDQ
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.236607 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.78 80 48.92 ;
    END
  END D_LVDS_I[2]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.558036 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.26 80 48.4 ;
    END
  END D_LVDS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_RTERMCAL_LVT28_H

MACRO RIIO_EG1D80V_RTERMCAL_RVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.46 80 40.6 ;
    END
  END VSSQ
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 567.2075 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 487.68 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 310.30352 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JV ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JW ;
    ANTENNAPARTIALCUTAREA 17.131488 LAYER A2 ;
    ANTENNADIFFAREA 152.2484 LAYER C4 ;
    ANTENNADIFFAREA 152.2484 LAYER C3 ;
    ANTENNADIFFAREA 152.2484 LAYER C5 ;
    ANTENNADIFFAREA 152.2484 LAYER JA ;
    ANTENNADIFFAREA 152.2484 LAYER QA ;
    ANTENNADIFFAREA 152.2484 LAYER QB ;
    ANTENNADIFFAREA 152.2484 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 98.217391 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.74 80 47.88 ;
    END
  END MODE_I[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 52.609456 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.22 80 47.36 ;
    END
  END MODE_I[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.7 80 46.84 ;
    END
  END RESULT_O[0]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.18 80 46.32 ;
    END
  END RESULT_O[1]
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.02 80 55.16 ;
    END
  END D_IOSG_I[10]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.811972 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.54 80 55.68 ;
    END
  END D_IOSG_I[11]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.82975 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.06 80 56.2 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C2 ;
      ANTENNAMAXAREACAR 14.865466 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.58 80 56.72 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C2 ;
      ANTENNAMAXAREACAR 14.455976 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.1 80 57.24 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C2 ;
      ANTENNAMAXAREACAR 13.688986 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.62 80 57.76 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.665245 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.34 80 50.48 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.666814 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.86 80 51 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.38 80 51.52 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.9 80 52.04 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.42 80 52.56 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.94 80 53.08 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.46 80 53.6 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.98 80 54.12 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 54.5 80 54.64 ;
    END
  END D_IOSG_I[9]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.629464 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.82 80 49.96 ;
    END
  END D_LVDS_I[0]
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.950893 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.3 80 49.44 ;
    END
  END D_LVDS_I[1]
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.98 80 41.12 ;
    END
  END VDDQ
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.236607 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.78 80 48.92 ;
    END
  END D_LVDS_I[2]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.558036 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.26 80 48.4 ;
    END
  END D_LVDS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_RTERMCAL_RVT28_H

MACRO RIIO_EG1D80V_RTERMCAL_SLVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_SLVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.46 80 40.6 ;
    END
  END VSSQ
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 567.2075 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 487.68 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 310.30352 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JV ;
    ANTENNAPARTIALCUTAREA 43.2 LAYER JW ;
    ANTENNAPARTIALCUTAREA 17.131488 LAYER A2 ;
    ANTENNADIFFAREA 152.2484 LAYER C4 ;
    ANTENNADIFFAREA 152.2484 LAYER C3 ;
    ANTENNADIFFAREA 152.2484 LAYER C5 ;
    ANTENNADIFFAREA 152.2484 LAYER JA ;
    ANTENNADIFFAREA 152.2484 LAYER QA ;
    ANTENNADIFFAREA 152.2484 LAYER QB ;
    ANTENNADIFFAREA 152.2484 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 98.217391 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.74 80 47.88 ;
    END
  END MODE_I[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 52.609456 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.22 80 47.36 ;
    END
  END MODE_I[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.7 80 46.84 ;
    END
  END RESULT_O[0]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.18 80 46.32 ;
    END
  END RESULT_O[1]
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.02 80 55.16 ;
    END
  END D_IOSG_I[10]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.811972 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.54 80 55.68 ;
    END
  END D_IOSG_I[11]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.82975 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.06 80 56.2 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C2 ;
      ANTENNAMAXAREACAR 14.865466 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.58 80 56.72 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C2 ;
      ANTENNAMAXAREACAR 14.455976 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.1 80 57.24 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C2 ;
      ANTENNAMAXAREACAR 13.688986 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.62 80 57.76 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.665245 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.34 80 50.48 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.666814 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.86 80 51 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.38 80 51.52 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.9 80 52.04 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.42 80 52.56 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.94 80 53.08 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.46 80 53.6 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.98 80 54.12 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 54.5 80 54.64 ;
    END
  END D_IOSG_I[9]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.629464 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.82 80 49.96 ;
    END
  END D_LVDS_I[0]
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.950893 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.3 80 49.44 ;
    END
  END D_LVDS_I[1]
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.98 80 41.12 ;
    END
  END VDDQ
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.236607 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.78 80 48.92 ;
    END
  END D_LVDS_I[2]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.558036 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.26 80 48.4 ;
    END
  END D_LVDS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_RTERMCAL_SLVT28_H

END LIBRARY
