----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 18.02.2022 13:47:38
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Noc_State_Machine_TB is
--  Port ( );
end Noc_State_Machine_TB;

architecture Behavioral of Noc_State_Machine_TB is
       
    component Noc_State_Machine
    port(
        clk                     : in  std_logic;
        Reset                   : in  std_logic;
        IO_data                 : in  std_logic_vector(127 downto 0);
        TAG_shift               : in  std_logic;                    
        TS                      : in  std_logic_vector(15 downto 0);
        PEC_Ready               : in  std_logic;
        Write_ack               : in  std_logic;
        FIFO_Ready1             : in  std_logic;
        FIFO_Ready2             : in  std_logic;
        FIFO_Ready3             : in  std_logic;        
        CMD_FF                  : in  std_logic;
        Opcode                  : in  std_logic_vector(11 downto 0);
        Loop_reg_mux_ctrl       : in  std_logic;        
        Load_RM_Address         : out std_logic;  
        Load_NOC_Reg            : out std_logic;  
        Load_PEC_Reg            : out std_logic;  
        Load_REQ_FF             : out std_logic; 
        En_IO_Data              : out std_logic;
        Load_GPP_CMD_Reg        : out std_logic;
        Reset_MDC               : out std_logic;
        Load_MD_Reg             : out std_logic;
        Step_MDC                : out std_logic;
        Sync_pulse              : out std_logic;
        En_RM                   : out std_logic;        
        Start_Tag_Shift         : out std_logic;                        
        Load_Tag_Shift_Counter  : out std_logic;                      
        Step_BC                 : out std_logic;  
        Reset_BC                : out std_logic;        
        Load_Mux_Reg            : out std_logic; 
        Control_Data_Out        : out std_logic_vector(7 downto 0);
        PEC_TS_Reg              : out std_logic_vector(15 downto 0);        
        Load_NOC_cmd_reg        : out std_logic;
        EN_TP_write             : out std_logic;
        EN_TP_read              : out std_logic;        
        Reset_TPC               : out std_logic;
        TP_Interchange          : out std_logic;
        En_IO_ctrl              : out std_logic;
        NOC_Ready               : out std_logic;
        load_Mode_reg           : out std_logic                              
      );
    end component;

    signal    clk                 : std_logic;
    signal    Reset               : std_logic;
    signal    IO_data             : std_logic_vector(127 downto 0);
    signal    TAG_shift           : std_logic;
    signal    TS                  : std_logic_vector(15 downto 0);
    signal    PEC_Ready           : std_logic;
    signal    Write_ack           : std_logic;
    signal    FIFO_ready1         : std_logic;
    signal    FIFO_ready2         : std_logic;
    signal    FIFO_ready3         : std_logic;
    signal    CMD_FF              : std_logic;
    signal    Opcode              : std_logic_vector(11 downto 0);
    signal    Loop_reg_mux_ctrl   : std_logic;
    signal    Load_RM_Address     : std_logic;
    signal    Load_NOC_Reg        : std_logic;
    signal    Load_PEC_Reg        : std_logic;
    signal    Load_REQ_FF         : std_logic;
    signal    En_IO_Data          : std_logic;
    signal    Load_GPP_CMD_Reg    : std_logic;
    signal    Reset_MDC           : std_logic;
    signal    Load_MD_Reg         : std_logic;
    signal    Step_MDC            : std_logic;
    signal    Sync_pulse          : std_logic;
    signal    En_RM               : std_logic;
    signal    Start_Tag_Shift     : std_logic;
    signal    Load_Tag_Shift_Counter  : std_logic;
    signal    Step_BC             : std_logic;
    signal    Reset_BC            : std_logic;
    signal    Load_Mux_Reg        : std_logic;
    signal    Control_Data_Out    : std_logic_vector(7 downto 0);
    signal    PEC_TS_Reg          : std_logic_vector(15 downto 0);        
    signal    Load_NOC_cmd_reg    : std_logic;
    signal    En_TP_write         : std_logic;
    signal    En_TP_read          : std_logic;
    signal    Reset_TPC           : std_logic;
    signal    TP_Interchange      : std_logic;
    signal    En_IO_ctrl          : std_logic;
    signal    NOC_Ready           : std_logic;
    signal    load_Mode_reg       : std_logic;
              
begin

    UUT: Noc_State_Machine port map (clk => clk, Reset => Reset, IO_data => IO_data, TAG_shift => TAG_shift, TS => TS, PEC_Ready => PEC_Ready, Write_ack => Write_ack, FIFO_ready1 => FIFO_ready1, FIFO_ready2 => FIFO_ready2, FIFO_ready3 => FIFO_ready3, CMD_FF => CMD_FF, Opcode => Opcode, Loop_reg_mux_ctrl => Loop_reg_mux_ctrl, Load_RM_Address => Load_RM_Address, Load_NOC_Reg => Load_NOC_Reg, Load_PEC_Reg => Load_PEC_Reg, Load_REQ_FF => Load_REQ_FF, En_IO_Data => En_IO_Data, Load_GPP_CMD_Reg => Load_GPP_CMD_Reg, Reset_MDC => Reset_MDC, Load_MD_Reg => Load_MD_Reg, Step_MDC => Step_MDC, Sync_pulse => Sync_pulse, En_RM => En_RM, Start_Tag_Shift => Start_Tag_Shift, Load_Tag_Shift_Counter => Load_Tag_Shift_Counter, Step_BC => Step_BC, Reset_BC => Reset_BC, Load_Mux_Reg => Load_Mux_Reg, Control_Data_Out => Control_Data_Out,  PEC_TS_Reg => PEC_TS_Reg, Load_NOC_cmd_reg => Load_NOC_cmd_reg, En_TP_write => En_TP_write, En_TP_read => En_TP_read, Reset_TPC => Reset_TPC, TP_Interchange => TP_Interchange, En_IO_ctrl => En_IO_ctrl, NOC_Ready => NOC_Ready, load_Mode_reg => load_Mode_reg);
 
    process
    begin
        Reset               <= '0';
        CMD_FF              <= '0';
        Write_ack           <= '0'; 
        FIFO_ready2         <= '0';
        fifo_ready3         <= '0';
        IO_data             <= (others => '0'); 
        Opcode              <= (others => '0');                                
        TS                  <= x"007D";
        TAG_shift           <= '0';
        Loop_reg_mux_ctrl   <= '0';  --comes from Mux reg
        wait for 50 ns;    
        Reset               <= '1';   
        wait for 40 ns;    
        Reset               <= '0';          
        wait for 300 ns;  
        CMD_FF              <= '1';           
        wait for 100 ns;
        CMD_FF              <= '0';  
        wait for 200 ns;
        Write_ack           <= '1';
        wait for 40 ns;
        Write_ack           <= '0';
        wait for 200 ns;
        FIFO_ready2         <= '1';
        wait for 100 ns;
        FIFO_ready2         <= '0';
        IO_data             <= x"00000000005000020000000000000000";
        wait for 100 ns;
        IO_data             <= x"0000070000C00203000C006000080001";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";      
        wait for 100 ns;
        IO_data             <= x"00080008001000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000660001000400000064800100040";  --40 is the address of command routine
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"08000608081000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000800062008100000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;        
        IO_data             <= x"00000000000000000000000000000000";       
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";          
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;        
        FIFO_ready2         <= '1';
        wait for 100 ns;
        FIFO_ready2         <= '0';
        IO_data             <= x"00000744081000F00000010200040012";  --81000f0 address write routine            
        wait for 100 ns;
        IO_data             <= x"000003080020000000000746081000E0"; --000003090020000000000746081000E0  LR=09 0r 08?
        wait for 100 ns;
        IO_data             <= x"00020000000000000250004900000103";
        wait for 100 ns;
        IO_data             <= x"04529055009E9004009E901400021000";
        wait for 100 ns;
        IO_data             <= x"000290000012904D000E902005529058";
        wait for 100 ns;
        IO_data             <= x"0000800000109049000E902000000000";  
        wait for 100 ns;
        IO_data             <= x"0000000000000000000480400010901A";   -- RM ->MUX-> DDR
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00020000000000000250006100000201";  
        wait for 100 ns;
        IO_data             <= x"0453D06D009FD004009FD01400035000"; 
        wait for 100 ns;
        IO_data             <= x"0003D2030013D965000FD0200553D070"; 
        wait for 100 ns;
        IO_data             <= x"000082030019D961000FD02000000000"; 
        wait for 100 ns;
        IO_data             <= x"009D9004000112030008030C0001D900"; 
        wait for 100 ns;
        IO_data             <= x"000000000004004000108000009D9004"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        -------------------------------------------------------------- 32 ta 0
        wait for 100 ns;        
        FIFO_ready2         <= '1';
        wait for 100 ns;
        FIFO_ready2         <= '0';
        IO_data             <= x"00000000000000000000000000000000";                 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;        
        FIFO_ready2         <= '1';
        wait for 100 ns;
        FIFO_ready2         <= '0';
        IO_data             <= x"00000000000000000000000000000000";                 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";                  
        --------------------------------------------------------------
        wait for 100 ns;        
        FIFO_ready2         <= '1';
        wait for 100 ns;
        FIFO_ready2         <= '0';
        IO_data             <= x"08000704081000F00000011100040012";  
        wait for 100 ns;
        IO_data             <= x"000003080020000008000706081000E0"; 
        wait for 100 ns;
        IO_data             <= x"0000800000008000000000000A500008"; 
        wait for 100 ns;
        IO_data             <= x"0C529015009E9004009E901400009000"; 
        wait for 100 ns;
        IO_data             <= x"0812900D00029000000E90200D52901A"; 
        wait for 100 ns;
        IO_data             <= x"0812100800021000000E902000029000"; 
        wait for 100 ns;
        IO_data             <= x"00121000000210000000000000020000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000060040"; 
        wait for 100 ns;         
        IO_data             <= x"00008000000000000A50002100000202";                 
        wait for 100 ns;
        IO_data             <= x"009FD004009FD0140000900000008000";
        wait for 100 ns;
        IO_data             <= x"000AD000000FD0200D5AD0350C5AD030";
        wait for 100 ns;
        IO_data             <= x"0000000000000000000AD203081AD026";
        wait for 100 ns;
        IO_data             <= x"081349210003500000035000000FD020";
        wait for 100 ns;
        IO_data             <= x"000349000003530D0003500000000203";  
        wait for 100 ns;
        IO_data             <= x"00100000009F0004009F000400000203";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000040040";  
        wait for 100 ns;
        FIFO_ready2         <= '1';
        wait for 100 ns;
        FIFO_ready2         <= '0';        
        IO_data             <= x"00000000000000000000000000000140";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000150"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;        
        IO_data             <= x"00000000000000000000000000000000";                 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        FIFO_ready2         <= '1';
        wait for 100 ns;
        FIFO_ready2         <= '0';        
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";                 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";        
        wait for 100 ns;
        FIFO_ready2         <= '1';
        wait for 100 ns;
        FIFO_ready2         <= '0';        
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";         
        wait for 100 ns;
        IO_data             <= x"0000000000000506081000E8000007F8"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000"; 
        wait for 100 ns;         
        IO_data             <= x"00000000000400300000000000040030";                 
        wait for 100 ns;
        IO_data             <= x"00000000003400300000000000040030";
        wait for 100 ns;
        IO_data             <= x"0030000000A0000000A0000000040001";
        wait for 100 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 100 ns;
        IO_data             <= x"0B5000F300080014000000000D5000F8";
        wait for 100 ns;
        IO_data             <= x"00000000000800040034000400000000";  
        wait for 100 ns;
        IO_data             <= x"00000000000000000004004000100000";                                                                                                                                                                                               
        wait for 200ns;
        CMD_FF              <= '1';
        Opcode              <= x"010";
        TS                  <= x"0010";    --Transfer size is 16 words            
        wait for 100 ns;
        CMD_FF              <= '0';
        wait for 160 ns;
        Write_ack           <= '1';
        wait for 100 ns;
        Write_ack           <= '0';
        -------------------------------------------------------------------------DATA IS READY IN FIFO
        wait for 380 ns;       
        FIFO_ready2         <= '1';
        wait for 80 ns;
        IO_data             <= x"00000000000000000000000000000000";
        wait for 20 ns;
        IO_data             <= x"11111111111111111111111111111111";        
        FIFO_ready2         <= '0';
        wait for 20 ns;
        IO_data             <= x"22222222222222222222222222222222";   
        wait for 20 ns;
        IO_data             <= x"33333333333333333333333333333333";
        wait for 20 ns;
        IO_data             <= x"44444444444444444444444444444444";
        wait for 20 ns;
        IO_data             <= x"55555555555555555555555555555555";        
        wait for 20 ns;
        IO_data             <= x"66666666666666666666666666666666";   
        wait for 20 ns;
        IO_data             <= x"77777777777777777777777777777777";
        wait for 20 ns;
        IO_data             <= x"88888888888888888888888888888888";
        wait for 20 ns;
        IO_data             <= x"99999999999999999999999999999999";        
        wait for 20 ns;
        IO_data             <= x"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";   
        wait for 20 ns;
        IO_data             <= x"BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB";
        wait for 20 ns;
        IO_data             <= x"CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC";
        wait for 20 ns;
        IO_data             <= x"DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD";        
        wait for 20 ns;
        IO_data             <= x"EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE";   
        wait for 20 ns;
        IO_data             <= x"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";                      
        wait for 200 ns;
        FIFO_ready3         <= '1';
        wait for 100 ns;
        FIFO_ready3         <= '0';
        wait for 220 ns;
        FIFO_ready3         <= '1';
        Write_ack           <= '1';
        wait for 100 ns;
        FIFO_ready3         <= '0';
        Write_ack           <= '0'; 
        wait for 220 ns;
        FIFO_ready3         <= '1';
        FIFO_ready2         <= '1';
        wait for 100 ns;
        FIFO_ready3         <= '0'; 
        wait for 220 ns;
        FIFO_ready3         <= '1';
        wait for 100 ns;
        FIFO_ready3         <= '0';
        wait for 220 ns;
        FIFO_ready3         <= '1';
        wait for 100 ns;
        FIFO_ready3         <= '0';
        wait for 220 ns;
        FIFO_ready3         <= '1';
        wait for 100 ns;
        FIFO_ready3         <= '0';
        wait for 220 ns;
        FIFO_ready3         <= '1';
        wait for 100 ns;
        FIFO_ready3         <= '0';                                                             
        wait for 1000000ns;           
    end process;
   
    process
    begin
        clk <= '0';
        for i in 1 to 100000 loop
            wait for 10ns;
            clk <= not clk;
        end loop;
        wait;
    end process;
    
end Behavioral;
