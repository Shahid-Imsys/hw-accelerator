use work.vetypes.all;
use work.instructiontypes.all;

entity ctrlmap_alu is
port (
  inst : in instruction;
  decoded : out all_addmul_ctrl);
end entity;

architecture generated of ctrlmap_alu is
begin
with inst select decoded <=
           (mux7l0 => L7, mux7l1 => L3, mux7r0 => onefft, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => zero, mux6r0 => onefft, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => L7, mux5l1 => L3, mux5r0 => onefft, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux4l0 => zero, mux4l1 => L2, mux4r0 => onefft, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L5, mux3l1 => L1, mux3r0 => onefft, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux1l0 => L5, mux1l1 => L1, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux0l0 => zero, mux0l1 => L0, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold)) when fftadd0,
           (mux7l0 => L7, mux7l1 => L3, mux7r0 => onefft, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux6l0 => L6, mux6l1 => zero, mux6r0 => onefft, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux5l0 => L7, mux5l1 => L3, mux5r0 => onefft, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux4l0 => zero, mux4l1 => L2, mux4r0 => onefft, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux3l0 => L5, mux3l1 => L1, mux3r0 => onefft, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L5, mux1l1 => L1, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux0l0 => zero, mux0l1 => L0, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable)) when fftadd1,
           (mux7l0 => L7, mux7l1 => L3, mux7r0 => R7, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => L2, mux6r0 => R7, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux5l0 => L7, mux5l1 => L3, mux5r0 => R6, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux4l0 => L6, mux4l1 => L2, mux4r0 => R6, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux3l0 => L5, mux3l1 => L1, mux3r0 => R5, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux2l0 => L4, mux2l1 => L0, mux2r0 => R5, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux1l0 => L5, mux1l1 => L1, mux1r0 => R4, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux0l0 => L4, mux0l1 => L0, mux0r0 => R4, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable)) when fftsub0,
           (mux7l0 => L7, mux7l1 => L3, mux7r0 => R5, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => L2, mux6r0 => R5, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux5l0 => L7, mux5l1 => L3, mux5r0 => R4, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux4l0 => L6, mux4l1 => L2, mux4r0 => R4, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux3l0 => L5, mux3l1 => L1, mux3r0 => R7, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux2l0 => L4, mux2l1 => L0, mux2r0 => R7, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux1l0 => L5, mux1l1 => L1, mux1r0 => R6, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux0l0 => L4, mux0l1 => L0, mux0r0 => R6, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable)) when fftsub1,
           (mux7l0 => L7, mux7l1 => ZpD, mux7r0 => R7, mux7r1 => ZpW,
            addmul7 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => ZpD, mux6r0 => R6, mux6r1 => ZpW,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux5l0 => L5, mux5l1 => ZpD, mux5r0 => R5, mux5r1 => ZpW,
            addmul5 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux4l0 => L4, mux4l1 => ZpD, mux4r0 => R4, mux4r1 => ZpW,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => ZpD, mux3r0 => R3, mux3r1 => ZpW,
            addmul3 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux2l0 => L2, mux2l1 => ZpD, mux2r0 => R2, mux2r1 => ZpW,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => ZpD, mux1r0 => R1, mux1r1 => ZpW,
            addmul1 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux0l0 => L0, mux0l1 => ZpD, mux0r0 => R0, mux0r1 => ZpW,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable)) when conv,
           (mux7l0 => L7, mux7l1 => ZpD, mux7r0 => R7, mux7r1 => ZpW,
            addmul7 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => ZpD, mux6r0 => R6, mux6r1 => ZpW,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux5l0 => L5, mux5l1 => ZpD, mux5r0 => R5, mux5r1 => ZpW,
            addmul5 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux4l0 => L4, mux4l1 => ZpD, mux4r0 => R4, mux4r1 => ZpW,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => ZpD, mux3r0 => R3, mux3r1 => ZpW,
            addmul3 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux2l0 => L2, mux2l1 => ZpD, mux2r0 => R2, mux2r1 => ZpW,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => ZpD, mux1r0 => R1, mux1r1 => ZpW,
            addmul1 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux0l0 => L0, mux0l1 => ZpD, mux0r0 => R0, mux0r1 => ZpW,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable)) when firstconv,
           (mux7l0 => L7, mux7l1 => ZpD, mux7r0 => R7, mux7r1 => ZpW,
            addmul7 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => ZpD, mux6r0 => R6, mux6r1 => ZpW,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux5l0 => L5, mux5l1 => ZpD, mux5r0 => R5, mux5r1 => ZpW,
            addmul5 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux4l0 => L4, mux4l1 => ZpD, mux4r0 => R4, mux4r1 => ZpW,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => ZpD, mux3r0 => R3, mux3r1 => ZpW,
            addmul3 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux2l0 => L2, mux2l1 => ZpD, mux2r0 => R2, mux2r1 => ZpW,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => ZpD, mux1r0 => R1, mux1r1 => ZpW,
            addmul1 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux0l0 => L0, mux0l1 => ZpD, mux0r0 => R0, mux0r1 => ZpW,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable)) when lastconv,
           (mux7l0 => L7, mux7l1 => ZpD, mux7r0 => R7, mux7r1 => ZpW,
            addmul7 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => ZpD, mux6r0 => R6, mux6r1 => ZpW,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux5l0 => L5, mux5l1 => ZpD, mux5r0 => R5, mux5r1 => ZpW,
            addmul5 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux4l0 => L4, mux4l1 => ZpD, mux4r0 => R4, mux4r1 => ZpW,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => ZpD, mux3r0 => R3, mux3r1 => ZpW,
            addmul3 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux2l0 => L2, mux2l1 => ZpD, mux2r0 => R2, mux2r1 => ZpW,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => ZpD, mux1r0 => R1, mux1r1 => ZpW,
            addmul1 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux0l0 => L0, mux0l1 => ZpD, mux0r0 => R0, mux0r1 => ZpW,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable)) when sum,
           (mux7l0 => L7, mux7l1 => ZpD, mux7r0 => R7, mux7r1 => ZpW,
            addmul7 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux6l0 => L6, mux6l1 => ZpD, mux6r0 => R6, mux6r1 => ZpW,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux5l0 => L5, mux5l1 => ZpD, mux5r0 => R5, mux5r1 => ZpW,
            addmul5 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux4l0 => L4, mux4l1 => ZpD, mux4r0 => R4, mux4r1 => ZpW,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux3l0 => L3, mux3l1 => ZpD, mux3r0 => R3, mux3r1 => ZpW,
            addmul3 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux2l0 => L2, mux2l1 => ZpD, mux2r0 => R2, mux2r1 => ZpW,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux1l0 => L1, mux1l1 => ZpD, mux1r0 => R1, mux1r1 => ZpW,
            addmul1 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux0l0 => L0, mux0l1 => ZpD, mux0r0 => R0, mux0r1 => ZpW,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold)) when nop,
           (mux7l0 => L7, mux7l1 => zero, mux7r0 => R7, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => zero, mux6r0 => R7, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => L7, mux5l1 => zero, mux5r0 => R6, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => L6, mux4l1 => zero, mux4r0 => R6, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L5, mux3l1 => zero, mux3r0 => R3, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => R3, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L5, mux1l1 => zero, mux1r0 => R2, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux0l0 => L4, mux0l1 => zero, mux0r0 => R2, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable)) when matmul00,
           (mux7l0 => L7, mux7l1 => zero, mux7r0 => R5, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => zero, mux6r0 => R5, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => L7, mux5l1 => zero, mux5r0 => R4, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => L6, mux4l1 => zero, mux4r0 => R4, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L5, mux3l1 => zero, mux3r0 => R1, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => R1, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L5, mux1l1 => zero, mux1r0 => R0, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux0l0 => L4, mux0l1 => zero, mux0r0 => R0, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable)) when matmul01,
           (mux7l0 => zero, mux7l1 => L3, mux7r0 => R5, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => zero, mux6l1 => L2, mux6r0 => R5, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => zero, mux5l1 => L3, mux5r0 => R4, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => zero, mux4l1 => L2, mux4r0 => R4, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => zero, mux3l1 => L1, mux3r0 => R1, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => zero, mux2l1 => L0, mux2r0 => R1, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => R0, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux0l0 => L0, mux0l1 => zero, mux0r0 => R0, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable)) when matmul11,
           (mux7l0 => zero, mux7l1 => L3, mux7r0 => R7, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => zero, mux6l1 => L2, mux6r0 => R7, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => zero, mux5l1 => L3, mux5r0 => R6, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => zero, mux4l1 => L2, mux4r0 => R6, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => zero, mux3l1 => L1, mux3r0 => R3, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => zero, mux2l1 => L0, mux2r0 => R3, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => R2, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux0l0 => L0, mux0l1 => zero, mux0r0 => R2, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable)) when matmul10,
           (mux7l0 => L7, mux7l1 => R7, mux7r0 => onefft, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => zero, mux6l1 => R6, mux6r0 => onefft, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => L5, mux5l1 => R5, mux5r0 => onefft, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux4l0 => L6, mux4l1 => zero, mux4r0 => onefft, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => R3, mux3r0 => onefft, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux1l0 => L1, mux1l1 => R1, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux0l0 => zero, mux0l1 => R0, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold)) when matadd00,
           (mux7l0 => L7, mux7l1 => R7, mux7r0 => onefft, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux6l0 => zero, mux6l1 => R6, mux6r0 => onefft, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux5l0 => L5, mux5l1 => R5, mux5r0 => onefft, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => zero, mux4l1 => R4, mux4r0 => onefft, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => R3, mux3r0 => onefft, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => R1, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux0l0 => zero, mux0l1 => R0, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold)) when matadd01,
           (mux7l0 => L7, mux7l1 => R7, mux7r0 => onefft, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux6l0 => zero, mux6l1 => R6, mux6r0 => onefft, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux5l0 => L5, mux5l1 => R5, mux5r0 => onefft, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux4l0 => zero, mux4l1 => L2, mux4r0 => onefft, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => R3, mux3r0 => onefft, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => zero, mux2l1 => R2, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => R1, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux0l0 => zero, mux0l1 => R0, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold)) when matadd10,
           (mux7l0 => L7, mux7l1 => R7, mux7r0 => onefft, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux6l0 => zero, mux6l1 => R6, mux6r0 => onefft, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux5l0 => L5, mux5l1 => R5, mux5r0 => onefft, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux4l0 => zero, mux4l1 => L2, mux4r0 => onefft, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux3l0 => L3, mux3l1 => R3, mux3r0 => onefft, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux2l0 => zero, mux2l1 => L0, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => R1, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux0l0 => zero, mux0l1 => R0, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable)) when matadd11,
           (mux7l0 => L7, mux7l1 => R7, mux7r0 => onefft, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => R6, mux6r0 => onefft, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux5l0 => L5, mux5l1 => R5, mux5r0 => onefft, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux4l0 => L4, mux4l1 => R4, mux4r0 => onefft, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => R3, mux3r0 => onefft, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux2l0 => L2, mux2l1 => R2, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => R1, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux0l0 => L0, mux0l1 => R0, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable)) when matsub,
           (mux7l0 => L7, mux7l1 => zero, mux7r0 => L1, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => zero, mux6r0 => L1, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => L7, mux5l1 => zero, mux5r0 => L0, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => L6, mux4l1 => zero, mux4r0 => L0, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux3l0 => L5, mux3l1 => zero, mux3r0 => L3, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => L3, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L5, mux1l1 => zero, mux1r0 => L2, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux0l0 => L4, mux0l1 => zero, mux0r0 => L2, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable)) when matdet,
           (mux7l0 => L7, mux7l1 => zero, mux7r0 => R7, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => zero, mux6r0 => R7, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => L7, mux5l1 => zero, mux5r0 => R6, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => L6, mux4l1 => zero, mux4r0 => R6, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L5, mux3l1 => zero, mux3r0 => R5, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => R5, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L5, mux1l1 => zero, mux1r0 => R4, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux0l0 => L4, mux0l1 => zero, mux0r0 => R4, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable)) when matmul00t,
           (mux7l0 => L7, mux7l1 => zero, mux7r0 => R3, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => zero, mux6r0 => R3, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => L7, mux5l1 => zero, mux5r0 => R2, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => L6, mux4l1 => zero, mux4r0 => R2, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L5, mux3l1 => zero, mux3r0 => R1, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => R1, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L5, mux1l1 => zero, mux1r0 => R0, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux0l0 => L4, mux0l1 => zero, mux0r0 => R0, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable)) when matmul01t,
           (mux7l0 => zero, mux7l1 => L3, mux7r0 => R3, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => zero, mux6l1 => L2, mux6r0 => R3, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => zero, mux5l1 => L3, mux5r0 => R2, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => zero, mux4l1 => L2, mux4r0 => R2, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => zero, mux3l1 => L1, mux3r0 => R1, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => zero, mux2l1 => L0, mux2r0 => R1, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => R0, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux0l0 => L0, mux0l1 => zero, mux0r0 => R0, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable)) when matmul11t,
           (mux7l0 => zero, mux7l1 => L3, mux7r0 => R7, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => zero, mux6l1 => L2, mux6r0 => R7, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => zero, mux5l1 => L3, mux5r0 => R6, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => zero, mux4l1 => L2, mux4r0 => R6, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => zero, mux3l1 => L1, mux3r0 => R5, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => zero, mux2l1 => L0, mux2r0 => R5, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => R4, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux0l0 => L0, mux0l1 => zero, mux0r0 => R4, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable)) when matmul10t,
           (mux7l0 => L7, mux7l1 => zero, mux7r0 => onefft, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => zero, mux6r0 => onefft, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U ,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => L7, mux5l1 => zero, mux5r0 => R2, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux4l0 => L6, mux4l1 => zero, mux4r0 => R2, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux3l0 => L5, mux3l1 => zero, mux3r0 => one, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => one, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux0l0 => zero, mux0l1 => zero, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold)) when unitri1,
           (mux7l0 => L7, mux7l1 => zero, mux7r0 => R3, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => L6, mux6l1 => zero, mux6r0 => R3, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => L7, mux5l1 => zero, mux5r0 => R2, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => L6, mux4l1 => zero, mux4r0 => R2, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L5, mux3l1 => zero, mux3r0 => one, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => L4, mux2l1 => zero, mux2r0 => one, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux0l0 => zero, mux0l1 => zero, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold)) when unitri2,
           (mux7l0 => zero, mux7l1 => L3, mux7r0 => onefft, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => zero, mux6l1 => L2, mux6r0 => onefft, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => zero, mux5l1 => L3, mux5r0 => R2, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux4l0 => zero, mux4l1 => L2, mux4r0 => R2, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux3l0 => zero, mux3l1 => L1, mux3r0 => one, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux2l0 => zero, mux2l1 => L0, mux2r0 => one, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux0l0 => zero, mux0l1 => zero, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold)) when unitri3,
           (mux7l0 => zero, mux7l1 => L3, mux7r0 => R3, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => zero, mux6l1 => L2, mux6r0 => R3, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => zero, mux5l1 => L3, mux5r0 => R2, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => zero, mux4l1 => L2, mux4r0 => R2, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => zero, mux3l1 => L1, mux3r0 => one, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => zero, mux2l1 => L0, mux2r0 => one, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux0l0 => zero, mux0l1 => zero, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold)) when unitri4,
            (mux7l0 => zero, mux7l1 => L5, mux7r0 => F3, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => zero, mux6l1 => L4, mux6r0 => F3, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => S, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => zero, mux5l1 => L5, mux5r0 => F2, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => zero, mux4l1 => L4, mux4r0 => F2, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => zero, mux3l1 => L1, mux3r0 => one, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => zero, mux2l1 => L0, mux2r0 => one, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux0l0 => zero, mux0l1 => zero, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold)) when unispec,
           (mux7l0 => L7, mux7l1 => zero, mux7r0 => onefft, mux7r1 => zero,
            addmul7 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable), -- TODO: add?
            mux6l0 => L6, mux6l1 => zero, mux6r0 => onefft, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux5l0 => L5, mux5l1 => zero, mux5r0 => onefft, mux5r1 => zero,
            addmul5 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux4l0 => L4, mux4l1 => zero, mux4r0 => onefft, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => zero, mux3r0 => onefft, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux2l0 => L2, mux2l1 => zero, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux0l0 => L0, mux0l1 => zero, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable)) when abs16,
           (mux7l0 => F7, mux7l1 => zero, mux7r0 => F1, mux7r1 => zero,
            addmul7 => (signl0 => U, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => F6, mux6l1 => zero, mux6r0 => F1, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => F7, mux5l1 => zero, mux5r0 => F0, mux5r1 => zero,
            addmul5 => (signl0 => U, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => F6, mux4l1 => zero, mux4r0 => F0, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => zero, mux3r0 => onefft, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux2l0 => L2, mux2l1 => zero, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux0l0 => L0, mux0l1 => zero, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold)) when mulden,
           (mux7l0 => F5, mux7l1 => zero, mux7r0 => F1, mux7r1 => zero,
            addmul7 => (signl0 => U, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => F4, mux6l1 => zero, mux6r0 => F1, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => F5, mux5l1 => zero, mux5r0 => F0, mux5r1 => zero,
            addmul5 => (signl0 => U, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => F4, mux4l1 => zero, mux4r0 => F0, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => L3, mux3l1 => zero, mux3r0 => onefft, mux3r1 => zero,
            addmul3 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => hold),
            mux2l0 => L2, mux2l1 => zero, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux0l0 => L0, mux0l1 => zero, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold)) when mulnum,
           (mux7l0 => F7, mux7l1 => zero, mux7r0 => F5, mux7r1 => zero,
            addmul7 => (signl0 => U, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux6l0 => F6, mux6l1 => zero, mux6r0 => F5, mux6r1 => zero,
            addmul6 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux5l0 => F7, mux5l1 => zero, mux5r0 => F4, mux5r1 => zero,
            addmul5 => (signl0 => U, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux4l0 => F6, mux4l1 => zero, mux4r0 => F4, mux4r1 => zero,
            addmul4 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux3l0 => F7, mux3l1 => zero, mux3r0 => onefft, mux3r1 => zero, --mux3r0 => x"02"
            addmul3 => (signl0 => U, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => add, addsubr => sub, en_addmul => enable),
            mux2l0 => F6, mux2l1 => zero, mux2r0 => onefft, mux2r1 => zero,
            addmul2 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => enable),
            mux1l0 => L1, mux1l1 => zero, mux1r0 => onefft, mux1r1 => zero,
            addmul1 => (signl0 => S, signl1 => S, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold),
            mux0l0 => L0, mux0l1 => zero, mux0r0 => onefft, mux0r1 => zero,
            addmul0 => (signl0 => U, signl1 => U, signr0 => U, signr1 => U,
                        addsubl => sub, addsubr => sub, en_addmul => hold)) when nrit;
end architecture;
