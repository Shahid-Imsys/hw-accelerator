VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


MACRO RIIO_EG1D80V_HPLVDS_RX_SLVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_HPLVDS_RX_SLVT28_V 0 0 ;
  SIZE 180 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN RTERM_TRIM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.348214 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.35 79.84 39.51 80 ;
    END
  END RTERM_TRIM_I[3]
  PIN RTERM_TRIM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.544643 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.71 79.84 35.87 80 ;
    END
  END RTERM_TRIM_I[2]
  PIN RTERM_TRIM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.741071 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 32.07 79.84 32.23 80 ;
    END
  END RTERM_TRIM_I[1]
  PIN RTERM_TRIM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.419643 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 28.43 79.84 28.59 80 ;
    END
  END RTERM_TRIM_I[0]
  PIN RTERM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.401664 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 27.91 79.84 28.07 80 ;
    END
  END RTERM_EN_I
  PIN RX_CTLE_RES_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8845 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1392 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 683.977778 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 93.43 79.84 93.59 80 ;
    END
  END RX_CTLE_RES_I[7]
  PIN RX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 64.31 79.84 64.47 80 ;
    END
  END RX_VCM_EN_I
  PIN DI_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNADIFFAREA 0.16192 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 67.43 79.84 67.59 80 ;
    END
  END DI_O
  PIN EI_DETECT_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 67.95 79.84 68.11 80 ;
    END
  END EI_DETECT_EN_I
  PIN RX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C1 ;
      ANTENNAMAXAREACAR 11.598214 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 69.51 79.84 69.67 80 ;
    END
  END RX_POL_I
  PIN RX_CTLE_CAP_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7795 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0336 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.256 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 872.669697 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 89.01 79.84 89.17 80 ;
    END
  END RX_CTLE_CAP_I[2]
  PIN RX_GAIN_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8215 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.208 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 385.255556 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 87.97 79.84 88.13 80 ;
    END
  END RX_GAIN_I[3]
  PIN RX_CTLE_RES_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8005 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0496 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.232 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 688.269697 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 91.35 79.84 91.51 80 ;
    END
  END RX_CTLE_RES_I[3]
  PIN RX_CTLE_RES_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8635 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1168 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 685.039394 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 92.91 79.84 93.07 80 ;
    END
  END RX_CTLE_RES_I[6]
  PIN RX_GAIN_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8635 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1168 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 385.923333 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 86.93 79.84 87.09 80 ;
    END
  END RX_GAIN_I[1]
  PIN RX_CTLE_RES_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7585 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0416 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 690.423232 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 90.31 79.84 90.47 80 ;
    END
  END RX_CTLE_RES_I[1]
  PIN RX_CTLE_CAP_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7585 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0416 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 896.394949 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 89.53 79.84 89.69 80 ;
    END
  END RX_CTLE_CAP_I[3]
  PIN RX_CTLE_RES_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7795 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.02744 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.256 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 689.346465 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 90.83 79.84 90.99 80 ;
    END
  END RX_CTLE_RES_I[2]
  PIN RX_GAIN_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0944 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.184 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 386.518889 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 87.45 79.84 87.61 80 ;
    END
  END RX_GAIN_I[2]
  PIN A_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3851.735 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 4546.871 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 2833.6725 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 3533.4 LAYER JA ;
    ANTENNAPARTIALMETALAREA 4709.88 LAYER OI ;
    ANTENNAPARTIALMETALAREA 35.36175 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 39.362752 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 38.123712 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 53.13276 LAYER YS ;
    ANTENNAPARTIALCUTAREA 84.610656 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.82224 LAYER A2 ;
    ANTENNADIFFAREA 889.8282 LAYER C4 ;
    ANTENNADIFFAREA 889.8282 LAYER C3 ;
    ANTENNADIFFAREA 889.8282 LAYER C5 ;
    ANTENNADIFFAREA 889.8282 LAYER JA ;
    ANTENNADIFFAREA 889.8282 LAYER OI ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    PORT
      LAYER C4 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
      LAYER JA ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 1.25 0 4.85 1.85 ;
      LAYER C5 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
      LAYER C2 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 1.25 0 4.85 1.85 ;
      LAYER OI ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 25.35 ;
        RECT 71.75 0 75.35 25.35 ;
        RECT 67.05 0 70.65 25.35 ;
        RECT 62.35 0 65.95 25.35 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 25.35 ;
        RECT 34.15 0 37.75 25.35 ;
        RECT 29.45 0 33.05 25.35 ;
        RECT 24.75 0 28.35 25.35 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 1.25 0 4.85 25.35 ;
      LAYER C3 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
    END
  END A_PAD_B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 10.95 78.15 13.95 80 ;
      LAYER OI ;
        RECT 10.95 78.15 13.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 15.65 78.15 18.65 80 ;
      LAYER OI ;
        RECT 15.65 78.15 18.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 29.75 78.15 32.75 80 ;
      LAYER OI ;
        RECT 29.75 78.15 32.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 34.45 78.15 37.45 80 ;
      LAYER OI ;
        RECT 34.45 78.15 37.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 48.55 78.15 51.55 80 ;
      LAYER OI ;
        RECT 48.55 78.15 51.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 53.25 78.15 56.25 80 ;
      LAYER OI ;
        RECT 53.25 78.15 56.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 67.35 78.15 70.35 80 ;
      LAYER OI ;
        RECT 67.35 78.15 70.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 72.05 78.15 75.05 80 ;
      LAYER OI ;
        RECT 72.05 78.15 75.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 86.15 78.15 89.15 80 ;
      LAYER OI ;
        RECT 86.15 78.15 89.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 90.85 78.15 93.85 80 ;
      LAYER OI ;
        RECT 90.85 78.15 93.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 104.95 78.15 107.95 80 ;
      LAYER OI ;
        RECT 104.95 78.15 107.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 109.65 78.15 112.65 80 ;
      LAYER OI ;
        RECT 109.65 78.15 112.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 123.75 78.15 126.75 80 ;
      LAYER OI ;
        RECT 123.75 78.15 126.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 128.45 78.15 131.45 80 ;
      LAYER OI ;
        RECT 128.45 78.15 131.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 142.55 78.15 145.55 80 ;
      LAYER OI ;
        RECT 142.55 78.15 145.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 147.25 78.15 150.25 80 ;
      LAYER OI ;
        RECT 147.25 78.15 150.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 161.35 78.15 164.35 80 ;
      LAYER OI ;
        RECT 161.35 78.15 164.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 166.05 78.15 169.05 80 ;
      LAYER OI ;
        RECT 166.05 78.15 169.05 80 ;
    END
    PORT
      LAYER JA ;
        RECT 0 68.75 180 72.35 ;
    END
    PORT
      LAYER JA ;
        RECT 0 64.05 180 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 1.55 78.15 4.55 80 ;
      LAYER OI ;
        RECT 1.55 78.15 4.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 6.25 78.15 9.25 80 ;
      LAYER OI ;
        RECT 6.25 78.15 9.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 20.35 78.15 23.35 80 ;
      LAYER OI ;
        RECT 20.35 78.15 23.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 25.05 78.15 28.05 80 ;
      LAYER OI ;
        RECT 25.05 78.15 28.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 39.15 78.15 42.15 80 ;
      LAYER OI ;
        RECT 39.15 78.15 42.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 43.85 78.15 46.85 80 ;
      LAYER OI ;
        RECT 43.85 78.15 46.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 57.95 78.15 60.95 80 ;
      LAYER OI ;
        RECT 57.95 78.15 60.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 62.65 78.15 65.65 80 ;
      LAYER OI ;
        RECT 62.65 78.15 65.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 76.75 78.15 79.75 80 ;
      LAYER OI ;
        RECT 76.75 78.15 79.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 81.45 78.15 84.45 80 ;
      LAYER OI ;
        RECT 81.45 78.15 84.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 95.55 78.15 98.55 80 ;
      LAYER OI ;
        RECT 95.55 78.15 98.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 100.25 78.15 103.25 80 ;
      LAYER OI ;
        RECT 100.25 78.15 103.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 114.35 78.15 117.35 80 ;
      LAYER OI ;
        RECT 114.35 78.15 117.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 119.05 78.15 122.05 80 ;
      LAYER OI ;
        RECT 119.05 78.15 122.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 133.15 78.15 136.15 80 ;
      LAYER OI ;
        RECT 133.15 78.15 136.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 137.85 78.15 140.85 80 ;
      LAYER OI ;
        RECT 137.85 78.15 140.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 151.95 78.15 154.95 80 ;
      LAYER OI ;
        RECT 151.95 78.15 154.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 156.65 78.15 159.65 80 ;
      LAYER OI ;
        RECT 156.65 78.15 159.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 170.75 78.15 173.75 80 ;
      LAYER OI ;
        RECT 170.75 78.15 173.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 175.45 78.15 178.45 80 ;
      LAYER OI ;
        RECT 175.45 78.15 178.45 80 ;
    END
    PORT
      LAYER JA ;
        RECT 0 73.45 180 77.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 59.35 180 62.95 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 0 54.65 180 58.25 ;
    END
    PORT
      LAYER JA ;
        RECT 0 45.25 180 48.85 ;
    END
    PORT
      LAYER JA ;
        RECT 0 40.55 180 44.15 ;
    END
    PORT
      LAYER JA ;
        RECT 0 26.45 180 30.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 17.05 180 20.65 ;
    END
    PORT
      LAYER JA ;
        RECT 0 3.67 180 6.55 ;
    END
  END VSSIO
  PIN B_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2385.0375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1287.3555 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 2651.475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 3059.37 LAYER JA ;
    ANTENNAPARTIALMETALAREA 3707.37 LAYER OI ;
    ANTENNAPARTIALMETALAREA 35.36175 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 24.45168 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.602784 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 170.367624 LAYER YS ;
    ANTENNAPARTIALCUTAREA 182.65824 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.82224 LAYER A2 ;
    ANTENNADIFFAREA 721.7962 LAYER C4 ;
    ANTENNADIFFAREA 334.12 LAYER C3 ;
    ANTENNADIFFAREA 721.7962 LAYER C5 ;
    ANTENNADIFFAREA 721.7962 LAYER JA ;
    ANTENNADIFFAREA 721.7962 LAYER OI ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    PORT
      LAYER C4 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER JA ;
        RECT 175.15 0 178.75 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C5 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C2 ;
        RECT 175.15 0 178.75 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER OI ;
        RECT 175.15 0 178.75 25.35 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 25.35 ;
        RECT 146.95 0 150.55 25.35 ;
        RECT 142.25 0 145.85 25.35 ;
        RECT 137.55 0 141.15 25.35 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 25.35 ;
        RECT 109.35 0 112.95 25.35 ;
        RECT 104.65 0 108.25 25.35 ;
        RECT 99.95 0 103.55 25.35 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C3 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
    END
  END B_PAD_B
  PIN RX_CTLE_CAP_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8005 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0496 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.232 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 873.912121 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 88.49 79.84 88.65 80 ;
    END
  END RX_CTLE_CAP_I[1]
  PIN RX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8845 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1392 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 384.76 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 86.41 79.84 86.57 80 ;
    END
  END RX_EN_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 0 49.95 180 53.55 ;
    END
    PORT
      LAYER JA ;
        RECT 0 35.85 180 39.45 ;
    END
    PORT
      LAYER JA ;
        RECT 0 31.15 180 34.75 ;
    END
    PORT
      LAYER JA ;
        RECT 0 12.35 180 15.95 ;
    END
    PORT
      LAYER JA ;
        RECT 0 7.65 180 11.25 ;
    END
  END VDDIO
  PIN EI_DETECT_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.01654 LAYER C1 ;
    ANTENNADIFFAREA 0.081 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 110.33 79.84 110.49 80 ;
    END
  END EI_DETECT_O
  PIN RX_CTLE_RES_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0944 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.184 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 686.116162 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 92.39 79.84 92.55 80 ;
    END
  END RX_CTLE_RES_I[5]
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.408 LAYER C4 ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER C4 ;
        RECT 0 39.575 180 40.825 ;
    END
  END VBIAS
  PIN RX_CTLE_RES_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8215 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.208 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 687.192929 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 91.87 79.84 92.03 80 ;
    END
  END RX_CTLE_RES_I[4]
  OBS
    LAYER CA ;
      RECT 0 0 180 80 ;
    LAYER M1 ;
      RECT 0 0 180 80 ;
    LAYER V1 ;
      RECT 0 0 180 80 ;
    LAYER M2 ;
      RECT 0 0 180 80 ;
    LAYER A1 ;
      RECT 0 0 180 80 ;
    LAYER C2 ;
      RECT 0 0 180 80 ;
    LAYER CB ;
      RECT 0 0 180 80 ;
    LAYER YS ;
      RECT 0 0 180 80 ;
    LAYER OI ;
      RECT 0 0 180 80 ;
    LAYER JQ ;
      RECT 0 0 180 80 ;
    LAYER JA ;
      RECT 0 0 180 80 ;
    LAYER AY ;
      RECT 0 0 180 80 ;
    LAYER C1 ;
      RECT 0 0 180 80 ;
    LAYER C5 ;
      RECT 0 0 180 80 ;
    LAYER C4 ;
      RECT 0 0 180 80 ;
    LAYER C3 ;
      RECT 0 0 180 80 ;
    LAYER A4 ;
      RECT 0 0 180 80 ;
    LAYER A3 ;
      RECT 0 0 180 80 ;
    LAYER A2 ;
      RECT 0 0 180 80 ;
  END
END RIIO_EG1D80V_HPLVDS_RX_SLVT28_V

MACRO RIIO_EG1D80V_HPLVDS_TX_SLVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_HPLVDS_TX_SLVT28_V 0 0 ;
  SIZE 180 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN RTERM_TRIM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.348214 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.35 79.84 39.51 80 ;
    END
  END RTERM_TRIM_I[3]
  PIN RTERM_TRIM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.544643 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.71 79.84 35.87 80 ;
    END
  END RTERM_TRIM_I[2]
  PIN RTERM_TRIM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.741071 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 32.07 79.84 32.23 80 ;
    END
  END RTERM_TRIM_I[1]
  PIN RTERM_TRIM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 45.419643 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 28.43 79.84 28.59 80 ;
    END
  END RTERM_TRIM_I[0]
  PIN RTERM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.401664 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 27.91 79.84 28.07 80 ;
    END
  END RTERM_EN_I
  PIN RX_CTLE_RES_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8845 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1392 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 683.977778 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 93.43 79.84 93.59 80 ;
    END
  END RX_CTLE_RES_I[7]
  PIN RX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 64.31 79.84 64.47 80 ;
    END
  END RX_VCM_EN_I
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C1 ;
      ANTENNAMAXAREACAR 11.288393 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.99 79.84 43.15 80 ;
    END
  END DO_I
  PIN DI_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNADIFFAREA 0.16192 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 67.43 79.84 67.59 80 ;
    END
  END DI_O
  PIN TX_BIAS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.446429 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 7.11 79.84 7.27 80 ;
    END
  END TX_BIAS_I[3]
  PIN EI_DETECT_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 67.95 79.84 68.11 80 ;
    END
  END EI_DETECT_EN_I
  PIN TX_BIAS_OD_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.23 79.84 23.39 80 ;
    END
  END TX_BIAS_OD_I
  PIN RX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C1 ;
      ANTENNAMAXAREACAR 11.598214 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 69.51 79.84 69.67 80 ;
    END
  END RX_POL_I
  PIN RX_CTLE_CAP_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7795 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0336 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.256 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 872.669697 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 89.01 79.84 89.17 80 ;
    END
  END RX_CTLE_CAP_I[2]
  PIN TX_VCM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.839286 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 55.47 79.84 55.63 80 ;
    END
  END TX_VCM_I[1]
  PIN RX_GAIN_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8215 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.208 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 385.255556 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 87.97 79.84 88.13 80 ;
    END
  END RX_GAIN_I[3]
  PIN RX_CTLE_RES_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8005 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0496 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.232 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 688.269697 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 91.35 79.84 91.51 80 ;
    END
  END RX_CTLE_RES_I[3]
  PIN RX_CTLE_RES_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8635 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1168 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 685.039394 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 92.91 79.84 93.07 80 ;
    END
  END RX_CTLE_RES_I[6]
  PIN RX_GAIN_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8635 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1168 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 385.923333 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 86.93 79.84 87.09 80 ;
    END
  END RX_GAIN_I[1]
  PIN RX_CTLE_RES_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7585 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0416 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 690.423232 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 90.31 79.84 90.47 80 ;
    END
  END RX_CTLE_RES_I[1]
  PIN TX_BIAS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.517857 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 18.03 79.84 18.19 80 ;
    END
  END TX_BIAS_I[0]
  PIN RX_CTLE_CAP_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7585 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0416 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 896.394949 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 89.53 79.84 89.69 80 ;
    END
  END RX_CTLE_CAP_I[3]
  PIN RX_CTLE_RES_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7795 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.02744 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.256 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 689.346465 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 90.83 79.84 90.99 80 ;
    END
  END RX_CTLE_RES_I[2]
  PIN RX_GAIN_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0944 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.184 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 386.518889 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 87.45 79.84 87.61 80 ;
    END
  END RX_GAIN_I[2]
  PIN A_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3851.735 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 4546.871 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 2833.6725 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 3533.4 LAYER JA ;
    ANTENNAPARTIALMETALAREA 4709.88 LAYER OI ;
    ANTENNAPARTIALMETALAREA 35.36175 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 39.362752 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 38.123712 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 53.13276 LAYER YS ;
    ANTENNAPARTIALCUTAREA 84.610656 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.82224 LAYER A2 ;
    ANTENNADIFFAREA 997.3482 LAYER C4 ;
    ANTENNADIFFAREA 997.3482 LAYER C3 ;
    ANTENNADIFFAREA 997.3482 LAYER C5 ;
    ANTENNADIFFAREA 997.3482 LAYER JA ;
    ANTENNADIFFAREA 997.3482 LAYER OI ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    PORT
      LAYER C4 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
      LAYER C5 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
      LAYER JA ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 1.25 0 4.85 1.85 ;
      LAYER C2 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 1.25 0 4.85 1.85 ;
      LAYER OI ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 25.35 ;
        RECT 71.75 0 75.35 25.35 ;
        RECT 67.05 0 70.65 25.35 ;
        RECT 62.35 0 65.95 25.35 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 25.35 ;
        RECT 34.15 0 37.75 25.35 ;
        RECT 29.45 0 33.05 25.35 ;
        RECT 24.75 0 28.35 25.35 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 1.25 0 4.85 25.35 ;
      LAYER C3 ;
        RECT 81.15 0 84.75 1.85 ;
        RECT 76.45 0 80.05 1.85 ;
        RECT 71.75 0 75.35 1.85 ;
        RECT 67.05 0 70.65 1.85 ;
        RECT 62.35 0 65.95 1.85 ;
        RECT 57.65 0 61.25 1.85 ;
        RECT 52.95 0 56.55 1.85 ;
        RECT 48.25 0 51.85 1.85 ;
        RECT 43.55 0 47.15 1.85 ;
        RECT 38.85 0 42.45 1.85 ;
        RECT 34.15 0 37.75 1.85 ;
        RECT 29.45 0 33.05 1.85 ;
        RECT 24.75 0 28.35 1.85 ;
        RECT 20.05 0 23.65 1.85 ;
        RECT 15.35 0 18.95 1.85 ;
        RECT 10.65 0 14.25 1.85 ;
        RECT 5.95 0 9.55 1.85 ;
        RECT 2.5 0 4.85 1.85 ;
    END
  END A_PAD_B
  PIN TX_BIAS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.642857 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.75 79.84 10.91 80 ;
    END
  END TX_BIAS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 10.95 78.15 13.95 80 ;
      LAYER OI ;
        RECT 10.95 78.15 13.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 15.65 78.15 18.65 80 ;
      LAYER OI ;
        RECT 15.65 78.15 18.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 29.75 78.15 32.75 80 ;
      LAYER OI ;
        RECT 29.75 78.15 32.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 34.45 78.15 37.45 80 ;
      LAYER OI ;
        RECT 34.45 78.15 37.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 48.55 78.15 51.55 80 ;
      LAYER OI ;
        RECT 48.55 78.15 51.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 53.25 78.15 56.25 80 ;
      LAYER OI ;
        RECT 53.25 78.15 56.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 67.35 78.15 70.35 80 ;
      LAYER OI ;
        RECT 67.35 78.15 70.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 72.05 78.15 75.05 80 ;
      LAYER OI ;
        RECT 72.05 78.15 75.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 86.15 78.15 89.15 80 ;
      LAYER OI ;
        RECT 86.15 78.15 89.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 90.85 78.15 93.85 80 ;
      LAYER OI ;
        RECT 90.85 78.15 93.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 104.95 78.15 107.95 80 ;
      LAYER OI ;
        RECT 104.95 78.15 107.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 109.65 78.15 112.65 80 ;
      LAYER OI ;
        RECT 109.65 78.15 112.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 123.75 78.15 126.75 80 ;
      LAYER OI ;
        RECT 123.75 78.15 126.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 128.45 78.15 131.45 80 ;
      LAYER OI ;
        RECT 128.45 78.15 131.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 142.55 78.15 145.55 80 ;
      LAYER OI ;
        RECT 142.55 78.15 145.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 147.25 78.15 150.25 80 ;
      LAYER OI ;
        RECT 147.25 78.15 150.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 161.35 78.15 164.35 80 ;
      LAYER OI ;
        RECT 161.35 78.15 164.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 166.05 78.15 169.05 80 ;
      LAYER OI ;
        RECT 166.05 78.15 169.05 80 ;
    END
    PORT
      LAYER JA ;
        RECT 0 68.75 180 72.35 ;
    END
    PORT
      LAYER JA ;
        RECT 0 64.05 180 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 1.55 78.15 4.55 80 ;
      LAYER OI ;
        RECT 1.55 78.15 4.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 6.25 78.15 9.25 80 ;
      LAYER OI ;
        RECT 6.25 78.15 9.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 20.35 78.15 23.35 80 ;
      LAYER OI ;
        RECT 20.35 78.15 23.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 25.05 78.15 28.05 80 ;
      LAYER OI ;
        RECT 25.05 78.15 28.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 39.15 78.15 42.15 80 ;
      LAYER OI ;
        RECT 39.15 78.15 42.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 43.85 78.15 46.85 80 ;
      LAYER OI ;
        RECT 43.85 78.15 46.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 57.95 78.15 60.95 80 ;
      LAYER OI ;
        RECT 57.95 78.15 60.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 62.65 78.15 65.65 80 ;
      LAYER OI ;
        RECT 62.65 78.15 65.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 76.75 78.15 79.75 80 ;
      LAYER OI ;
        RECT 76.75 78.15 79.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 81.45 78.15 84.45 80 ;
      LAYER OI ;
        RECT 81.45 78.15 84.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 95.55 78.15 98.55 80 ;
      LAYER OI ;
        RECT 95.55 78.15 98.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 100.25 78.15 103.25 80 ;
      LAYER OI ;
        RECT 100.25 78.15 103.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 114.35 78.15 117.35 80 ;
      LAYER OI ;
        RECT 114.35 78.15 117.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 119.05 78.15 122.05 80 ;
      LAYER OI ;
        RECT 119.05 78.15 122.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 133.15 78.15 136.15 80 ;
      LAYER OI ;
        RECT 133.15 78.15 136.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 137.85 78.15 140.85 80 ;
      LAYER OI ;
        RECT 137.85 78.15 140.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 151.95 78.15 154.95 80 ;
      LAYER OI ;
        RECT 151.95 78.15 154.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 156.65 78.15 159.65 80 ;
      LAYER OI ;
        RECT 156.65 78.15 159.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 170.75 78.15 173.75 80 ;
      LAYER OI ;
        RECT 170.75 78.15 173.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 175.45 78.15 178.45 80 ;
      LAYER OI ;
        RECT 175.45 78.15 178.45 80 ;
    END
    PORT
      LAYER JA ;
        RECT 0 73.45 180 77.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 59.35 180 62.95 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 0 54.65 180 58.25 ;
    END
    PORT
      LAYER JA ;
        RECT 0 45.25 180 48.85 ;
    END
    PORT
      LAYER JA ;
        RECT 0 40.55 180 44.15 ;
    END
    PORT
      LAYER JA ;
        RECT 0 26.45 180 30.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 17.05 180 20.65 ;
    END
    PORT
      LAYER JA ;
        RECT 0 3.67 180 6.55 ;
    END
  END VSSIO
  PIN B_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2385.0375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1287.3555 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 2651.475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 3059.37 LAYER JA ;
    ANTENNAPARTIALMETALAREA 3707.37 LAYER OI ;
    ANTENNAPARTIALMETALAREA 35.36175 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 24.45168 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.602784 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 170.367624 LAYER YS ;
    ANTENNAPARTIALCUTAREA 182.65824 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.82224 LAYER A2 ;
    ANTENNADIFFAREA 775.5562 LAYER C4 ;
    ANTENNADIFFAREA 387.88 LAYER C3 ;
    ANTENNADIFFAREA 775.5562 LAYER C5 ;
    ANTENNADIFFAREA 775.5562 LAYER JA ;
    ANTENNADIFFAREA 775.5562 LAYER OI ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    PORT
      LAYER C4 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C5 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER JA ;
        RECT 175.15 0 178.75 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C2 ;
        RECT 175.15 0 178.75 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER OI ;
        RECT 175.15 0 178.75 25.35 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 25.35 ;
        RECT 146.95 0 150.55 25.35 ;
        RECT 142.25 0 145.85 25.35 ;
        RECT 137.55 0 141.15 25.35 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 25.35 ;
        RECT 109.35 0 112.95 25.35 ;
        RECT 104.65 0 108.25 25.35 ;
        RECT 99.95 0 103.55 25.35 ;
        RECT 95.25 0 98.85 1.85 ;
      LAYER C3 ;
        RECT 175.15 0 177.5 1.85 ;
        RECT 170.45 0 174.05 1.85 ;
        RECT 165.75 0 169.35 1.85 ;
        RECT 161.05 0 164.65 1.85 ;
        RECT 156.35 0 159.95 1.85 ;
        RECT 151.65 0 155.25 1.85 ;
        RECT 146.95 0 150.55 1.85 ;
        RECT 142.25 0 145.85 1.85 ;
        RECT 137.55 0 141.15 1.85 ;
        RECT 132.85 0 136.45 1.85 ;
        RECT 128.15 0 131.75 1.85 ;
        RECT 123.45 0 127.05 1.85 ;
        RECT 118.75 0 122.35 1.85 ;
        RECT 114.05 0 117.65 1.85 ;
        RECT 109.35 0 112.95 1.85 ;
        RECT 104.65 0 108.25 1.85 ;
        RECT 99.95 0 103.55 1.85 ;
        RECT 95.25 0 98.85 1.85 ;
    END
  END B_PAD_B
  PIN RX_CTLE_CAP_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8005 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0496 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.232 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 873.912121 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 88.49 79.84 88.65 80 ;
    END
  END RX_CTLE_CAP_I[1]
  PIN RX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8845 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.1392 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C3 ;
      ANTENNAMAXAREACAR 384.76 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 86.41 79.84 86.57 80 ;
    END
  END RX_EN_I
  PIN TX_VCM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.517857 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 59.11 79.84 59.27 80 ;
    END
  END TX_VCM_I[0]
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 0 49.95 180 53.55 ;
    END
    PORT
      LAYER JA ;
        RECT 0 35.85 180 39.45 ;
    END
    PORT
      LAYER JA ;
        RECT 0 31.15 180 34.75 ;
    END
    PORT
      LAYER JA ;
        RECT 0 12.35 180 15.95 ;
    END
    PORT
      LAYER JA ;
        RECT 0 7.65 180 11.25 ;
    END
  END VDDIO
  PIN TX_BIAS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.839286 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.39 79.84 14.55 80 ;
    END
  END TX_BIAS_I[1]
  PIN EI_DETECT_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.01654 LAYER C1 ;
    ANTENNADIFFAREA 0.081 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 110.33 79.84 110.49 80 ;
    END
  END EI_DETECT_O
  PIN TX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C1 ;
      ANTENNAMAXAREACAR 12.119643 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.47 79.84 42.63 80 ;
    END
  END TX_POL_I
  PIN RX_CTLE_RES_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.0944 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.184 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 686.116162 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 92.39 79.84 92.55 80 ;
    END
  END RX_CTLE_RES_I[5]
  PIN TX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.304261 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 60.67 79.84 60.83 80 ;
    END
  END TX_VCM_EN_I
  PIN RX_CTLE_RES_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8215 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 0.072 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 0.208 LAYER C1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.00396 LAYER A2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C3 ;
      ANTENNAMAXAREACAR 687.192929 LAYER C3 ;
    PORT
      LAYER C1 ;
        RECT 91.87 79.84 92.03 80 ;
    END
  END RX_CTLE_RES_I[4]
  PIN TX_VCM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.446429 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 48.19 79.84 48.35 80 ;
    END
  END TX_VCM_I[3]
  PIN TX_VCM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.642857 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 51.83 79.84 51.99 80 ;
    END
  END TX_VCM_I[2]
  PIN TX_EI_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0112 LAYER C1 ;
      ANTENNAMAXAREACAR 22.714286 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 45.33 79.84 45.49 80 ;
    END
  END TX_EI_I
  PIN TX_FFE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2048 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02128 LAYER C1 ;
      ANTENNAMAXAREACAR 14.671992 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 49.23 79.84 49.39 80 ;
    END
  END TX_FFE_I
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.408 LAYER C4 ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER C4 ;
        RECT 0 39.575 180 40.825 ;
    END
  END VBIAS
  PIN TX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.304261 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.59 79.84 19.75 80 ;
    END
  END TX_EN_I
  OBS
    LAYER CA ;
      RECT 0 0 180 80 ;
    LAYER M1 ;
      RECT 0 0 180 80 ;
    LAYER V1 ;
      RECT 0 0 180 80 ;
    LAYER M2 ;
      RECT 0 0 180 80 ;
    LAYER A1 ;
      RECT 0 0 180 80 ;
    LAYER C2 ;
      RECT 0 0 180 80 ;
    LAYER CB ;
      RECT 0 0 180 80 ;
    LAYER YS ;
      RECT 0 0 180 80 ;
    LAYER OI ;
      RECT 0 0 180 80 ;
    LAYER JQ ;
      RECT 0 0 180 80 ;
    LAYER JA ;
      RECT 0 0 180 80 ;
    LAYER AY ;
      RECT 0 0 180 80 ;
    LAYER C1 ;
      RECT 0 0 180 80 ;
    LAYER C5 ;
      RECT 0 0 180 80 ;
    LAYER C4 ;
      RECT 0 0 180 80 ;
    LAYER C3 ;
      RECT 0 0 180 80 ;
    LAYER A4 ;
      RECT 0 0 180 80 ;
    LAYER A3 ;
      RECT 0 0 180 80 ;
    LAYER A2 ;
      RECT 0 0 180 80 ;
  END
END RIIO_EG1D80V_HPLVDS_TX_SLVT28_V

MACRO RIIO_EG1D80V_RTERMCAL_HVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_HVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 59.35 60 62.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER JA ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER JA ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER JA ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER JA ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER JA ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER JA ;
        RECT 54.35 78.15 57.35 80 ;
    END
  END VSS
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.564137 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.2 79.86 40.34 80 ;
    END
  END D_IOSG_I[10]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2212 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.36 79.86 5.5 80 ;
    END
  END RESULT_O[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.84 79.86 4.98 80 ;
    END
  END RESULT_O[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.336729 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.4 79.86 19.54 80 ;
    END
  END MODE_I[1]
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.869565 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.04 79.86 23.18 80 ;
    END
  END MODE_I[0]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.058036 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.92 79.86 7.06 80 ;
    END
  END D_LVDS_I[3]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER JA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER JA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER JA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER JA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.736607 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.56 79.86 10.7 80 ;
    END
  END D_LVDS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER JA ;
        RECT 0 64.05 60 67.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER JA ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER JA ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER JA ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER JA ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER JA ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER JA ;
        RECT 49.65 78.15 52.65 80 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER JA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER JA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER JA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER JA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 68.1725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 389.395 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER JA ;
    ANTENNAPARTIALMETALAREA 603.245 LAYER OI ;
    ANTENNAPARTIALMETALAREA 235.02 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.5176 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 26.737776 LAYER YS ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 7.031552 LAYER A2 ;
    ANTENNADIFFAREA 167.0608 LAYER C4 ;
    ANTENNADIFFAREA 167.0608 LAYER C3 ;
    ANTENNADIFFAREA 167.0608 LAYER C5 ;
    ANTENNADIFFAREA 167.0608 LAYER JA ;
    ANTENNADIFFAREA 167.0608 LAYER OI ;
    ANTENNADIFFAREA 167.0608 LAYER C2 ;
    PORT
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.84 79.86 30.98 80 ;
    END
  END VDDQ
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.450893 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.2 79.86 14.34 80 ;
    END
  END D_LVDS_I[1]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.129464 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.84 79.86 17.98 80 ;
    END
  END D_LVDS_I[0]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.637946 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.68 79.86 39.82 80 ;
    END
  END D_IOSG_I[9]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.518659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.16 79.86 39.3 80 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.594022 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.64 79.86 38.78 80 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.369792 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.12 79.86 38.26 80 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.446458 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.6 79.86 37.74 80 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.136806 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.08 79.86 37.22 80 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.214583 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.56 79.86 36.7 80 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.670735 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.04 79.86 36.18 80 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.747794 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.52 79.86 35.66 80 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C1 ;
      ANTENNAMAXAREACAR 2.443131 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.8 79.86 42.94 80 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C1 ;
      ANTENNAMAXAREACAR 2.582738 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.28 79.86 42.42 80 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C1 ;
      ANTENNAMAXAREACAR 2.733211 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.76 79.86 41.9 80 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.179861 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.24 79.86 41.38 80 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.253194 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.72 79.86 40.86 80 ;
    END
  END D_IOSG_I[11]
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.32 79.86 30.46 80 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_RTERMCAL_HVT28_V

MACRO RIIO_EG1D80V_RTERMCAL_LLHVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_LLHVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 59.35 60 62.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER JA ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER JA ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER JA ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER JA ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER JA ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER JA ;
        RECT 54.35 78.15 57.35 80 ;
    END
  END VSS
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.564137 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.2 79.86 40.34 80 ;
    END
  END D_IOSG_I[10]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2212 LAYER C1 ;
    ANTENNADIFFAREA 0.03864 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.36 79.86 5.5 80 ;
    END
  END RESULT_O[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNADIFFAREA 0.03864 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.84 79.86 4.98 80 ;
    END
  END RESULT_O[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.044 LAYER C1 ;
      ANTENNAMAXAREACAR 22.719659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.4 79.86 19.54 80 ;
    END
  END MODE_I[1]
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0184 LAYER C1 ;
      ANTENNAMAXAREACAR 19.954348 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.04 79.86 23.18 80 ;
    END
  END MODE_I[0]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C1 ;
      ANTENNAMAXAREACAR 59.65625 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.92 79.86 7.06 80 ;
    END
  END D_LVDS_I[3]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER JA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER JA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER JA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER JA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C1 ;
      ANTENNAMAXAREACAR 59.65625 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.56 79.86 10.7 80 ;
    END
  END D_LVDS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER JA ;
        RECT 0 64.05 60 67.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER JA ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER JA ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER JA ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER JA ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER JA ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER JA ;
        RECT 49.65 78.15 52.65 80 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER JA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER JA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER JA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER JA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 68.1725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 389.395 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER JA ;
    ANTENNAPARTIALMETALAREA 603.245 LAYER OI ;
    ANTENNAPARTIALMETALAREA 235.02 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.5176 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 26.737776 LAYER YS ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 7.031552 LAYER A2 ;
    ANTENNADIFFAREA 167.0608 LAYER C4 ;
    ANTENNADIFFAREA 167.0608 LAYER C3 ;
    ANTENNADIFFAREA 167.0608 LAYER C5 ;
    ANTENNADIFFAREA 167.0608 LAYER JA ;
    ANTENNADIFFAREA 167.0608 LAYER OI ;
    ANTENNADIFFAREA 167.0608 LAYER C2 ;
    PORT
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.84 79.86 30.98 80 ;
    END
  END VDDQ
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C1 ;
      ANTENNAMAXAREACAR 59.65625 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.2 79.86 14.34 80 ;
    END
  END D_LVDS_I[1]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C1 ;
      ANTENNAMAXAREACAR 60.30625 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.84 79.86 17.98 80 ;
    END
  END D_LVDS_I[0]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.637946 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.68 79.86 39.82 80 ;
    END
  END D_IOSG_I[9]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.518659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.16 79.86 39.3 80 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.594022 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.64 79.86 38.78 80 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.369792 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.12 79.86 38.26 80 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.446458 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.6 79.86 37.74 80 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.136806 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.08 79.86 37.22 80 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.214583 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.56 79.86 36.7 80 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.670735 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.04 79.86 36.18 80 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.747794 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.52 79.86 35.66 80 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C1 ;
      ANTENNAMAXAREACAR 2.443131 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.8 79.86 42.94 80 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C1 ;
      ANTENNAMAXAREACAR 2.582738 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.28 79.86 42.42 80 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C1 ;
      ANTENNAMAXAREACAR 2.733211 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.76 79.86 41.9 80 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.179861 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.24 79.86 41.38 80 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.253194 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.72 79.86 40.86 80 ;
    END
  END D_IOSG_I[11]
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.32 79.86 30.46 80 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_RTERMCAL_LLHVT28_V

MACRO RIIO_EG1D80V_RTERMCAL_LVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_LVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 59.35 60 62.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER JA ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER JA ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER JA ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER JA ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER JA ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER JA ;
        RECT 54.35 78.15 57.35 80 ;
    END
  END VSS
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.564137 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.2 79.86 40.34 80 ;
    END
  END D_IOSG_I[10]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2212 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.36 79.86 5.5 80 ;
    END
  END RESULT_O[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.84 79.86 4.98 80 ;
    END
  END RESULT_O[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.336729 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.4 79.86 19.54 80 ;
    END
  END MODE_I[1]
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.869565 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.04 79.86 23.18 80 ;
    END
  END MODE_I[0]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.058036 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.92 79.86 7.06 80 ;
    END
  END D_LVDS_I[3]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER JA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER JA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER JA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER JA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.736607 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.56 79.86 10.7 80 ;
    END
  END D_LVDS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER JA ;
        RECT 0 64.05 60 67.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER JA ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER JA ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER JA ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER JA ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER JA ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER JA ;
        RECT 49.65 78.15 52.65 80 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER JA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER JA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER JA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER JA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 68.1725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 389.395 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER JA ;
    ANTENNAPARTIALMETALAREA 603.245 LAYER OI ;
    ANTENNAPARTIALMETALAREA 235.02 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.5176 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 26.737776 LAYER YS ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 7.031552 LAYER A2 ;
    ANTENNADIFFAREA 167.0608 LAYER C4 ;
    ANTENNADIFFAREA 167.0608 LAYER C3 ;
    ANTENNADIFFAREA 167.0608 LAYER C5 ;
    ANTENNADIFFAREA 167.0608 LAYER JA ;
    ANTENNADIFFAREA 167.0608 LAYER OI ;
    ANTENNADIFFAREA 167.0608 LAYER C2 ;
    PORT
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.84 79.86 30.98 80 ;
    END
  END VDDQ
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.450893 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.2 79.86 14.34 80 ;
    END
  END D_LVDS_I[1]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.129464 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.84 79.86 17.98 80 ;
    END
  END D_LVDS_I[0]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.637946 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.68 79.86 39.82 80 ;
    END
  END D_IOSG_I[9]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.518659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.16 79.86 39.3 80 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.594022 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.64 79.86 38.78 80 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.369792 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.12 79.86 38.26 80 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.446458 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.6 79.86 37.74 80 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.136806 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.08 79.86 37.22 80 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.214583 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.56 79.86 36.7 80 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.670735 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.04 79.86 36.18 80 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.747794 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.52 79.86 35.66 80 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C1 ;
      ANTENNAMAXAREACAR 2.443131 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.8 79.86 42.94 80 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C1 ;
      ANTENNAMAXAREACAR 2.582738 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.28 79.86 42.42 80 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C1 ;
      ANTENNAMAXAREACAR 2.733211 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.76 79.86 41.9 80 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.179861 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.24 79.86 41.38 80 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.253194 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.72 79.86 40.86 80 ;
    END
  END D_IOSG_I[11]
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.32 79.86 30.46 80 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_RTERMCAL_LVT28_V

MACRO RIIO_EG1D80V_RTERMCAL_RVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 59.35 60 62.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER JA ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER JA ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER JA ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER JA ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER JA ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER JA ;
        RECT 54.35 78.15 57.35 80 ;
    END
  END VSS
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.564137 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.2 79.86 40.34 80 ;
    END
  END D_IOSG_I[10]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2212 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.36 79.86 5.5 80 ;
    END
  END RESULT_O[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.84 79.86 4.98 80 ;
    END
  END RESULT_O[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.336729 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.4 79.86 19.54 80 ;
    END
  END MODE_I[1]
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.869565 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.04 79.86 23.18 80 ;
    END
  END MODE_I[0]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.058036 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.92 79.86 7.06 80 ;
    END
  END D_LVDS_I[3]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER JA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER JA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER JA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER JA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.736607 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.56 79.86 10.7 80 ;
    END
  END D_LVDS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER JA ;
        RECT 0 64.05 60 67.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER JA ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER JA ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER JA ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER JA ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER JA ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER JA ;
        RECT 49.65 78.15 52.65 80 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER JA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER JA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER JA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER JA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 68.1725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 389.395 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER JA ;
    ANTENNAPARTIALMETALAREA 603.245 LAYER OI ;
    ANTENNAPARTIALMETALAREA 235.02 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.5176 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 26.737776 LAYER YS ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 7.031552 LAYER A2 ;
    ANTENNADIFFAREA 167.0608 LAYER C4 ;
    ANTENNADIFFAREA 167.0608 LAYER C3 ;
    ANTENNADIFFAREA 167.0608 LAYER C5 ;
    ANTENNADIFFAREA 167.0608 LAYER JA ;
    ANTENNADIFFAREA 167.0608 LAYER OI ;
    ANTENNADIFFAREA 167.0608 LAYER C2 ;
    PORT
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.84 79.86 30.98 80 ;
    END
  END VDDQ
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.450893 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.2 79.86 14.34 80 ;
    END
  END D_LVDS_I[1]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.129464 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.84 79.86 17.98 80 ;
    END
  END D_LVDS_I[0]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.637946 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.68 79.86 39.82 80 ;
    END
  END D_IOSG_I[9]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.518659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.16 79.86 39.3 80 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.594022 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.64 79.86 38.78 80 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.369792 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.12 79.86 38.26 80 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.446458 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.6 79.86 37.74 80 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.136806 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.08 79.86 37.22 80 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.214583 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.56 79.86 36.7 80 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.670735 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.04 79.86 36.18 80 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.747794 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.52 79.86 35.66 80 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C1 ;
      ANTENNAMAXAREACAR 2.443131 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.8 79.86 42.94 80 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C1 ;
      ANTENNAMAXAREACAR 2.582738 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.28 79.86 42.42 80 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C1 ;
      ANTENNAMAXAREACAR 2.733211 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.76 79.86 41.9 80 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.179861 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.24 79.86 41.38 80 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.253194 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.72 79.86 40.86 80 ;
    END
  END D_IOSG_I[11]
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.32 79.86 30.46 80 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_RTERMCAL_RVT28_V

MACRO RIIO_EG1D80V_RTERMCAL_SLVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_SLVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 59.35 60 62.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER JA ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER JA ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER JA ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER JA ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER JA ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER JA ;
        RECT 54.35 78.15 57.35 80 ;
    END
  END VSS
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.564137 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.2 79.86 40.34 80 ;
    END
  END D_IOSG_I[10]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2212 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.36 79.86 5.5 80 ;
    END
  END RESULT_O[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 4.84 79.86 4.98 80 ;
    END
  END RESULT_O[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C1 ;
      ANTENNAMAXAREACAR 17.336729 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.4 79.86 19.54 80 ;
    END
  END MODE_I[1]
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 13.869565 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.04 79.86 23.18 80 ;
    END
  END MODE_I[0]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.058036 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.92 79.86 7.06 80 ;
    END
  END D_LVDS_I[3]
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER JA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER JA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER JA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER JA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER JA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 43.736607 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.56 79.86 10.7 80 ;
    END
  END D_LVDS_I[2]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER JA ;
        RECT 0 64.05 60 67.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER JA ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER JA ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER JA ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER JA ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER JA ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER JA ;
        RECT 49.65 78.15 52.65 80 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER JA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER JA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER JA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER JA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 68.1725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 389.395 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER JA ;
    ANTENNAPARTIALMETALAREA 603.245 LAYER OI ;
    ANTENNAPARTIALMETALAREA 235.02 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 5.5176 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 26.737776 LAYER YS ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 7.031552 LAYER A2 ;
    ANTENNADIFFAREA 167.0608 LAYER C4 ;
    ANTENNADIFFAREA 167.0608 LAYER C3 ;
    ANTENNADIFFAREA 167.0608 LAYER C5 ;
    ANTENNADIFFAREA 167.0608 LAYER JA ;
    ANTENNADIFFAREA 167.0608 LAYER OI ;
    ANTENNADIFFAREA 167.0608 LAYER C2 ;
    PORT
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.84 79.86 30.98 80 ;
    END
  END VDDQ
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.450893 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.2 79.86 14.34 80 ;
    END
  END D_LVDS_I[1]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.322 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C1 ;
      ANTENNAMAXAREACAR 44.129464 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.84 79.86 17.98 80 ;
    END
  END D_LVDS_I[0]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C1 ;
      ANTENNAMAXAREACAR 3.637946 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.68 79.86 39.82 80 ;
    END
  END D_IOSG_I[9]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.518659 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.16 79.86 39.3 80 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C1 ;
      ANTENNAMAXAREACAR 4.594022 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.64 79.86 38.78 80 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.369792 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.12 79.86 38.26 80 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C1 ;
      ANTENNAMAXAREACAR 5.446458 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.6 79.86 37.74 80 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.136806 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.08 79.86 37.22 80 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C1 ;
      ANTENNAMAXAREACAR 6.214583 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.56 79.86 36.7 80 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.670735 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 36.04 79.86 36.18 80 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C1 ;
      ANTENNAMAXAREACAR 6.747794 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 35.52 79.86 35.66 80 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C1 ;
      ANTENNAMAXAREACAR 2.443131 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.8 79.86 42.94 80 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C1 ;
      ANTENNAMAXAREACAR 2.582738 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 42.28 79.86 42.42 80 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C1 ;
      ANTENNAMAXAREACAR 2.733211 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.76 79.86 41.9 80 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.179861 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 41.24 79.86 41.38 80 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51058 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C1 ;
      ANTENNAMAXAREACAR 3.253194 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.72 79.86 40.86 80 ;
    END
  END D_IOSG_I[11]
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 30.32 79.86 30.46 80 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_RTERMCAL_SLVT28_V


MACRO RIIO_EG1D80V_HPLVDS_RX_SLVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_HPLVDS_RX_SLVT28_H 0 0 ;
  SIZE 80 BY 180 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN A_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1022.5375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1004.7775 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 155.5575 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 467.37 LAYER JA ;
    ANTENNAPARTIALMETALAREA 36.63 LAYER OI ;
    ANTENNAPARTIALMETALAREA 748.6275 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 19.085088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 17.86928 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 6.170256 LAYER YS ;
    ANTENNAPARTIALCUTAREA 40.520736 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.713824 LAYER A2 ;
    ANTENNADIFFAREA 153.2196 LAYER C4 ;
    ANTENNADIFFAREA 153.2196 LAYER C3 ;
    ANTENNADIFFAREA 153.2196 LAYER C5 ;
    ANTENNADIFFAREA 153.2196 LAYER JA ;
    ANTENNADIFFAREA 153.2196 LAYER OI ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER C3 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER C4 ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 99.95 1.85 103.55 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER C5 ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 99.95 1.85 103.55 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER JA ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 99.95 1.85 103.55 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 178.75 ;
      LAYER OI ;
        RECT 0 99.95 25.35 103.55 ;
        RECT 0 104.65 25.35 108.25 ;
        RECT 0 109.35 25.35 112.95 ;
        RECT 0 114.05 25.35 117.65 ;
        RECT 0 137.55 25.35 141.15 ;
        RECT 0 142.25 25.35 145.85 ;
        RECT 0 146.95 25.35 150.55 ;
        RECT 0 151.65 25.35 155.25 ;
        RECT 0 175.15 25.35 178.75 ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
    END
  END A_PAD_B
  PIN RX_CTLE_RES_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7195 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.639394 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 91.09 80 91.25 ;
    END
  END RX_CTLE_RES_I[2]
  PIN RX_CTLE_RES_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6755 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.756566 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 90.57 80 90.73 ;
    END
  END RX_CTLE_RES_I[1]
  PIN RX_CTLE_RES_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9395 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 473.457576 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 93.69 80 93.85 ;
    END
  END RX_CTLE_RES_I[7]
  PIN RX_CTLE_CAP_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7635 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 468.536364 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 88.23 80 88.39 ;
    END
  END RX_CTLE_CAP_I[1]
  PIN RX_CTLE_CAP_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6755 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 478.89798 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 89.27 80 89.43 ;
    END
  END RX_CTLE_CAP_I[3]
  PIN RX_GAIN_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8515 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 347.915 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 87.19 80 87.35 ;
    END
  END RX_GAIN_I[2]
  PIN RX_CTLE_CAP_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7195 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 463.455556 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 88.75 80 88.91 ;
    END
  END RX_CTLE_CAP_I[2]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 59.35 0 62.95 180 ;
    END
    PORT
      LAYER JA ;
        RECT 73.45 0 77.05 180 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 175.45 80 178.45 ;
      LAYER OI ;
        RECT 78.15 175.45 80 178.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 170.75 80 173.75 ;
      LAYER OI ;
        RECT 78.15 170.75 80 173.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 156.65 80 159.65 ;
      LAYER OI ;
        RECT 78.15 156.65 80 159.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 151.95 80 154.95 ;
      LAYER OI ;
        RECT 78.15 151.95 80 154.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 137.85 80 140.85 ;
      LAYER OI ;
        RECT 78.15 137.85 80 140.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 133.15 80 136.15 ;
      LAYER OI ;
        RECT 78.15 133.15 80 136.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 119.05 80 122.05 ;
      LAYER OI ;
        RECT 78.15 119.05 80 122.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 114.35 80 117.35 ;
      LAYER OI ;
        RECT 78.15 114.35 80 117.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 100.25 80 103.25 ;
      LAYER OI ;
        RECT 78.15 100.25 80 103.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 95.55 80 98.55 ;
      LAYER OI ;
        RECT 78.15 95.55 80 98.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 81.45 80 84.45 ;
      LAYER OI ;
        RECT 78.15 81.45 80 84.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 76.75 80 79.75 ;
      LAYER OI ;
        RECT 78.15 76.75 80 79.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 62.65 80 65.65 ;
      LAYER OI ;
        RECT 78.15 62.65 80 65.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 57.95 80 60.95 ;
      LAYER OI ;
        RECT 78.15 57.95 80 60.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 43.85 80 46.85 ;
      LAYER OI ;
        RECT 78.15 43.85 80 46.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 39.15 80 42.15 ;
      LAYER OI ;
        RECT 78.15 39.15 80 42.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 25.05 80 28.05 ;
      LAYER OI ;
        RECT 78.15 25.05 80 28.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 20.35 80 23.35 ;
      LAYER OI ;
        RECT 78.15 20.35 80 23.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 6.25 80 9.25 ;
      LAYER OI ;
        RECT 78.15 6.25 80 9.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 1.55 80 4.55 ;
      LAYER OI ;
        RECT 78.15 1.55 80 4.55 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.408 LAYER C4 ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER C4 ;
        RECT 39.575 0 40.825 180 ;
    END
  END VBIAS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 3.67 0 6.55 180 ;
    END
    PORT
      LAYER JA ;
        RECT 17.05 0 20.65 180 ;
    END
    PORT
      LAYER JA ;
        RECT 26.45 0 30.05 180 ;
    END
    PORT
      LAYER JA ;
        RECT 40.55 0 44.15 180 ;
    END
    PORT
      LAYER JA ;
        RECT 45.25 0 48.85 180 ;
    END
    PORT
      LAYER JA ;
        RECT 54.65 0 58.25 180 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 7.65 0 11.25 180 ;
    END
    PORT
      LAYER JA ;
        RECT 12.35 0 15.95 180 ;
    END
    PORT
      LAYER JA ;
        RECT 31.15 0 34.75 180 ;
    END
    PORT
      LAYER JA ;
        RECT 35.85 0 39.45 180 ;
    END
    PORT
      LAYER JA ;
        RECT 49.95 0 53.55 180 ;
    END
  END VDDIO
  PIN RX_CTLE_RES_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8955 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 471.867677 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 93.17 80 93.33 ;
    END
  END RX_CTLE_RES_I[6]
  PIN RX_GAIN_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8955 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 347.558333 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 86.67 80 86.83 ;
    END
  END RX_GAIN_I[1]
  PIN EI_DETECT_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 35.102484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 131.91 80 132.07 ;
    END
  END EI_DETECT_EN_I
  PIN B_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1022.5375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1004.7775 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1090.5675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 467.37 LAYER JA ;
    ANTENNAPARTIALMETALAREA 826.65 LAYER OI ;
    ANTENNAPARTIALMETALAREA 747.92 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 19.085088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 17.86928 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 38.735496 LAYER YS ;
    ANTENNAPARTIALCUTAREA 41.570496 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.713824 LAYER A2 ;
    ANTENNADIFFAREA 153.2196 LAYER C4 ;
    ANTENNADIFFAREA 153.2196 LAYER C3 ;
    ANTENNADIFFAREA 153.2196 LAYER C5 ;
    ANTENNADIFFAREA 153.2196 LAYER JA ;
    ANTENNADIFFAREA 153.2196 LAYER OI ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
      LAYER C3 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
      LAYER C4 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
        RECT 0 76.45 1.85 80.05 ;
        RECT 0 81.15 1.85 84.75 ;
      LAYER C5 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
        RECT 0 76.45 1.85 80.05 ;
        RECT 0 81.15 1.85 84.75 ;
      LAYER JA ;
        RECT 0 1.25 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
        RECT 0 76.45 1.85 80.05 ;
        RECT 0 81.15 1.85 84.75 ;
      LAYER OI ;
        RECT 0 1.25 25.35 4.85 ;
        RECT 0 24.75 25.35 28.35 ;
        RECT 0 29.45 25.35 33.05 ;
        RECT 0 34.15 25.35 37.75 ;
        RECT 0 38.85 25.35 42.45 ;
        RECT 0 62.35 25.35 65.95 ;
        RECT 0 67.05 25.35 70.65 ;
        RECT 0 71.75 25.35 75.35 ;
        RECT 0 76.45 25.35 80.05 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 81.15 1.85 84.75 ;
    END
  END B_PAD_B
  PIN RX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 35.102484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 132.95 80 133.11 ;
    END
  END RX_VCM_EN_I
  PIN RX_CTLE_RES_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8515 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.287879 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 92.65 80 92.81 ;
    END
  END RX_CTLE_RES_I[5]
  PIN RX_CTLE_RES_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7635 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.522222 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 91.61 80 91.77 ;
    END
  END RX_CTLE_RES_I[3]
  PIN RX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9395 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 346.633889 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 86.15 80 86.31 ;
    END
  END RX_EN_I
  PIN RX_GAIN_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8075 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 346.412778 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 87.71 80 87.87 ;
    END
  END RX_GAIN_I[3]
  PIN DI_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2128 LAYER C2 ;
    ANTENNADIFFAREA 0.16192 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 129.83 80 129.99 ;
    END
  END DI_O
  PIN EI_DETECT_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2128 LAYER C2 ;
    ANTENNADIFFAREA 0.081 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 49.23 80 49.39 ;
    END
  END EI_DETECT_O
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 64.05 0 67.65 180 ;
    END
    PORT
      LAYER JA ;
        RECT 68.75 0 72.35 180 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 166.05 80 169.05 ;
      LAYER OI ;
        RECT 78.15 166.05 80 169.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 161.35 80 164.35 ;
      LAYER OI ;
        RECT 78.15 161.35 80 164.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 147.25 80 150.25 ;
      LAYER OI ;
        RECT 78.15 147.25 80 150.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 142.55 80 145.55 ;
      LAYER OI ;
        RECT 78.15 142.55 80 145.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 128.45 80 131.45 ;
      LAYER OI ;
        RECT 78.15 128.45 80 131.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 123.75 80 126.75 ;
      LAYER OI ;
        RECT 78.15 123.75 80 126.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 109.65 80 112.65 ;
      LAYER OI ;
        RECT 78.15 109.65 80 112.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 104.95 80 107.95 ;
      LAYER OI ;
        RECT 78.15 104.95 80 107.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 90.85 80 93.85 ;
      LAYER OI ;
        RECT 78.15 90.85 80 93.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 86.15 80 89.15 ;
      LAYER OI ;
        RECT 78.15 86.15 80 89.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 72.05 80 75.05 ;
      LAYER OI ;
        RECT 78.15 72.05 80 75.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 67.35 80 70.35 ;
      LAYER OI ;
        RECT 78.15 67.35 80 70.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 53.25 80 56.25 ;
      LAYER OI ;
        RECT 78.15 53.25 80 56.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 48.55 80 51.55 ;
      LAYER OI ;
        RECT 78.15 48.55 80 51.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 34.45 80 37.45 ;
      LAYER OI ;
        RECT 78.15 34.45 80 37.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 29.75 80 32.75 ;
      LAYER OI ;
        RECT 78.15 29.75 80 32.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 15.65 80 18.65 ;
      LAYER OI ;
        RECT 78.15 15.65 80 18.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 10.95 80 13.95 ;
      LAYER OI ;
        RECT 78.15 10.95 80 13.95 ;
    END
  END VDD
  PIN RX_CTLE_RES_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8075 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.405051 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 92.13 80 92.29 ;
    END
  END RX_CTLE_RES_I[4]
  PIN RTERM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 28.891274 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 175.07 80 175.23 ;
    END
  END RTERM_EN_I
  PIN RTERM_TRIM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 175.59 80 175.75 ;
    END
  END RTERM_TRIM_I[0]
  PIN RTERM_TRIM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 176.11 80 176.27 ;
    END
  END RTERM_TRIM_I[1]
  PIN RTERM_TRIM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 176.63 80 176.79 ;
    END
  END RTERM_TRIM_I[2]
  PIN RTERM_TRIM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 177.15 80 177.31 ;
    END
  END RTERM_TRIM_I[3]
  PIN RX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C2 ;
      ANTENNAMAXAREACAR 56.869643 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 128.27 80 128.43 ;
    END
  END RX_POL_I
  OBS
    LAYER CA ;
      RECT 0 0 80 180 ;
    LAYER M1 ;
      RECT 0 0 80 180 ;
    LAYER V1 ;
      RECT 0 0 80 180 ;
    LAYER M2 ;
      RECT 0 0 80 180 ;
    LAYER A1 ;
      RECT 0 0 80 180 ;
    LAYER C2 ;
      RECT 0 0 80 180 ;
    LAYER CB ;
      RECT 0 0 80 180 ;
    LAYER YS ;
      RECT 0 0 80 180 ;
    LAYER OI ;
      RECT 0 0 80 180 ;
    LAYER JQ ;
      RECT 0 0 80 180 ;
    LAYER JA ;
      RECT 0 0 80 180 ;
    LAYER AY ;
      RECT 0 0 80 180 ;
    LAYER C1 ;
      RECT 0 0 80 180 ;
    LAYER C5 ;
      RECT 0 0 80 180 ;
    LAYER C4 ;
      RECT 0 0 80 180 ;
    LAYER C3 ;
      RECT 0 0 80 180 ;
    LAYER A4 ;
      RECT 0 0 80 180 ;
    LAYER A3 ;
      RECT 0 0 80 180 ;
    LAYER A2 ;
      RECT 0 0 80 180 ;
  END
END RIIO_EG1D80V_HPLVDS_RX_SLVT28_H

MACRO RIIO_EG1D80V_HPLVDS_TX_SLVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_HPLVDS_TX_SLVT28_H 0 0 ;
  SIZE 80 BY 180 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN A_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1022.5375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1004.7775 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 155.5575 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 467.37 LAYER JA ;
    ANTENNAPARTIALMETALAREA 36.63 LAYER OI ;
    ANTENNAPARTIALMETALAREA 748.6275 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 19.085088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 17.86928 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 6.170256 LAYER YS ;
    ANTENNAPARTIALCUTAREA 40.520736 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.713824 LAYER A2 ;
    ANTENNADIFFAREA 206.9796 LAYER C4 ;
    ANTENNADIFFAREA 206.9796 LAYER C3 ;
    ANTENNADIFFAREA 206.9796 LAYER C5 ;
    ANTENNADIFFAREA 206.9796 LAYER JA ;
    ANTENNADIFFAREA 206.9796 LAYER OI ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER C3 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER C4 ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 99.95 1.85 103.55 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER C5 ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 99.95 1.85 103.55 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 177.5 ;
      LAYER JA ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 99.95 1.85 103.55 ;
        RECT 0 104.65 1.85 108.25 ;
        RECT 0 109.35 1.85 112.95 ;
        RECT 0 114.05 1.85 117.65 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 137.55 1.85 141.15 ;
        RECT 0 142.25 1.85 145.85 ;
        RECT 0 146.95 1.85 150.55 ;
        RECT 0 151.65 1.85 155.25 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
        RECT 0 175.15 1.85 178.75 ;
      LAYER OI ;
        RECT 0 99.95 25.35 103.55 ;
        RECT 0 104.65 25.35 108.25 ;
        RECT 0 109.35 25.35 112.95 ;
        RECT 0 114.05 25.35 117.65 ;
        RECT 0 137.55 25.35 141.15 ;
        RECT 0 142.25 25.35 145.85 ;
        RECT 0 146.95 25.35 150.55 ;
        RECT 0 151.65 25.35 155.25 ;
        RECT 0 175.15 25.35 178.75 ;
        RECT 0 95.25 1.85 98.85 ;
        RECT 0 118.75 1.85 122.35 ;
        RECT 0 123.45 1.85 127.05 ;
        RECT 0 128.15 1.85 131.75 ;
        RECT 0 132.85 1.85 136.45 ;
        RECT 0 156.35 1.85 159.95 ;
        RECT 0 161.05 1.85 164.65 ;
        RECT 0 165.75 1.85 169.35 ;
        RECT 0 170.45 1.85 174.05 ;
    END
  END A_PAD_B
  PIN RX_CTLE_RES_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7195 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.639394 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 91.09 80 91.25 ;
    END
  END RX_CTLE_RES_I[2]
  PIN RX_CTLE_RES_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6755 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.756566 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 90.57 80 90.73 ;
    END
  END RX_CTLE_RES_I[1]
  PIN RX_CTLE_RES_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9395 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 473.457576 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 93.69 80 93.85 ;
    END
  END RX_CTLE_RES_I[7]
  PIN TX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 32.20556 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 148.55 80 148.71 ;
    END
  END TX_VCM_EN_I
  PIN RX_CTLE_CAP_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7635 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 468.536364 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 88.23 80 88.39 ;
    END
  END RX_CTLE_CAP_I[1]
  PIN RX_CTLE_CAP_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6755 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 478.89798 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 89.27 80 89.43 ;
    END
  END RX_CTLE_CAP_I[3]
  PIN TX_BIAS_OD_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 35.102484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 132.43 80 132.59 ;
    END
  END TX_BIAS_OD_I
  PIN RX_GAIN_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8515 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 347.915 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 87.19 80 87.35 ;
    END
  END RX_GAIN_I[2]
  PIN RX_CTLE_CAP_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7195 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 463.455556 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 88.75 80 88.91 ;
    END
  END RX_CTLE_CAP_I[2]
  PIN TX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C2 ;
      ANTENNAMAXAREACAR 54.698214 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 127.75 80 127.91 ;
    END
  END TX_POL_I
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 59.35 0 62.95 180 ;
    END
    PORT
      LAYER JA ;
        RECT 73.45 0 77.05 180 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 175.45 80 178.45 ;
      LAYER OI ;
        RECT 78.15 175.45 80 178.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 170.75 80 173.75 ;
      LAYER OI ;
        RECT 78.15 170.75 80 173.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 156.65 80 159.65 ;
      LAYER OI ;
        RECT 78.15 156.65 80 159.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 151.95 80 154.95 ;
      LAYER OI ;
        RECT 78.15 151.95 80 154.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 137.85 80 140.85 ;
      LAYER OI ;
        RECT 78.15 137.85 80 140.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 133.15 80 136.15 ;
      LAYER OI ;
        RECT 78.15 133.15 80 136.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 119.05 80 122.05 ;
      LAYER OI ;
        RECT 78.15 119.05 80 122.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 114.35 80 117.35 ;
      LAYER OI ;
        RECT 78.15 114.35 80 117.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 100.25 80 103.25 ;
      LAYER OI ;
        RECT 78.15 100.25 80 103.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 95.55 80 98.55 ;
      LAYER OI ;
        RECT 78.15 95.55 80 98.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 81.45 80 84.45 ;
      LAYER OI ;
        RECT 78.15 81.45 80 84.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 76.75 80 79.75 ;
      LAYER OI ;
        RECT 78.15 76.75 80 79.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 62.65 80 65.65 ;
      LAYER OI ;
        RECT 78.15 62.65 80 65.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 57.95 80 60.95 ;
      LAYER OI ;
        RECT 78.15 57.95 80 60.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 43.85 80 46.85 ;
      LAYER OI ;
        RECT 78.15 43.85 80 46.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 39.15 80 42.15 ;
      LAYER OI ;
        RECT 78.15 39.15 80 42.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 25.05 80 28.05 ;
      LAYER OI ;
        RECT 78.15 25.05 80 28.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 20.35 80 23.35 ;
      LAYER OI ;
        RECT 78.15 20.35 80 23.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 6.25 80 9.25 ;
      LAYER OI ;
        RECT 78.15 6.25 80 9.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 1.55 80 4.55 ;
      LAYER OI ;
        RECT 78.15 1.55 80 4.55 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.408 LAYER C4 ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER C4 ;
        RECT 39.575 0 40.825 180 ;
    END
  END VBIAS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 3.67 0 6.55 180 ;
    END
    PORT
      LAYER JA ;
        RECT 17.05 0 20.65 180 ;
    END
    PORT
      LAYER JA ;
        RECT 26.45 0 30.05 180 ;
    END
    PORT
      LAYER JA ;
        RECT 40.55 0 44.15 180 ;
    END
    PORT
      LAYER JA ;
        RECT 45.25 0 48.85 180 ;
    END
    PORT
      LAYER JA ;
        RECT 54.65 0 58.25 180 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 7.65 0 11.25 180 ;
    END
    PORT
      LAYER JA ;
        RECT 12.35 0 15.95 180 ;
    END
    PORT
      LAYER JA ;
        RECT 31.15 0 34.75 180 ;
    END
    PORT
      LAYER JA ;
        RECT 35.85 0 39.45 180 ;
    END
    PORT
      LAYER JA ;
        RECT 49.95 0 53.55 180 ;
    END
  END VDDIO
  PIN RX_CTLE_RES_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8955 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 471.867677 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 93.17 80 93.33 ;
    END
  END RX_CTLE_RES_I[6]
  PIN RX_GAIN_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8955 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 347.558333 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 86.67 80 86.83 ;
    END
  END RX_GAIN_I[1]
  PIN TX_BIAS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 152.71 80 152.87 ;
    END
  END TX_BIAS_I[2]
  PIN TX_VCM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 149.07 80 149.23 ;
    END
  END TX_VCM_I[0]
  PIN EI_DETECT_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 35.102484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 131.91 80 132.07 ;
    END
  END EI_DETECT_EN_I
  PIN B_PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1022.5375 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1004.7775 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1090.5675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 467.37 LAYER JA ;
    ANTENNAPARTIALMETALAREA 826.65 LAYER OI ;
    ANTENNAPARTIALMETALAREA 747.92 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 19.085088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 17.86928 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 38.735496 LAYER YS ;
    ANTENNAPARTIALCUTAREA 41.570496 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.713824 LAYER A2 ;
    ANTENNADIFFAREA 206.9796 LAYER C4 ;
    ANTENNADIFFAREA 206.9796 LAYER C3 ;
    ANTENNADIFFAREA 206.9796 LAYER C5 ;
    ANTENNADIFFAREA 206.9796 LAYER JA ;
    ANTENNADIFFAREA 206.9796 LAYER OI ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
      LAYER C3 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
      LAYER C4 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
        RECT 0 76.45 1.85 80.05 ;
        RECT 0 81.15 1.85 84.75 ;
      LAYER C5 ;
        RECT 0 2.5 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
        RECT 0 76.45 1.85 80.05 ;
        RECT 0 81.15 1.85 84.75 ;
      LAYER JA ;
        RECT 0 1.25 1.85 4.85 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 24.75 1.85 28.35 ;
        RECT 0 29.45 1.85 33.05 ;
        RECT 0 34.15 1.85 37.75 ;
        RECT 0 38.85 1.85 42.45 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 62.35 1.85 65.95 ;
        RECT 0 67.05 1.85 70.65 ;
        RECT 0 71.75 1.85 75.35 ;
        RECT 0 76.45 1.85 80.05 ;
        RECT 0 81.15 1.85 84.75 ;
      LAYER OI ;
        RECT 0 1.25 25.35 4.85 ;
        RECT 0 24.75 25.35 28.35 ;
        RECT 0 29.45 25.35 33.05 ;
        RECT 0 34.15 25.35 37.75 ;
        RECT 0 38.85 25.35 42.45 ;
        RECT 0 62.35 25.35 65.95 ;
        RECT 0 67.05 25.35 70.65 ;
        RECT 0 71.75 25.35 75.35 ;
        RECT 0 76.45 25.35 80.05 ;
        RECT 0 5.95 1.85 9.55 ;
        RECT 0 10.65 1.85 14.25 ;
        RECT 0 15.35 1.85 18.95 ;
        RECT 0 20.05 1.85 23.65 ;
        RECT 0 43.55 1.85 47.15 ;
        RECT 0 48.25 1.85 51.85 ;
        RECT 0 52.95 1.85 56.55 ;
        RECT 0 57.65 1.85 61.25 ;
        RECT 0 81.15 1.85 84.75 ;
    END
  END B_PAD_B
  PIN RX_VCM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 35.102484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 132.95 80 133.11 ;
    END
  END RX_VCM_EN_I
  PIN TX_VCM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 149.59 80 149.75 ;
    END
  END TX_VCM_I[1]
  PIN RX_CTLE_RES_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8515 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.287879 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 92.65 80 92.81 ;
    END
  END RX_CTLE_RES_I[5]
  PIN TX_VCM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 150.63 80 150.79 ;
    END
  END TX_VCM_I[3]
  PIN RX_CTLE_RES_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7635 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.522222 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 91.61 80 91.77 ;
    END
  END RX_CTLE_RES_I[3]
  PIN RX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9395 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 346.633889 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 86.15 80 86.31 ;
    END
  END RX_EN_I
  PIN TX_VCM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 150.11 80 150.27 ;
    END
  END TX_VCM_I[2]
  PIN TX_EI_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0112 LAYER C2 ;
      ANTENNAMAXAREACAR 99.871429 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 128.79 80 128.95 ;
    END
  END TX_EI_I
  PIN TX_BIAS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 151.67 80 151.83 ;
    END
  END TX_BIAS_I[0]
  PIN TX_BIAS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 152.19 80 152.35 ;
    END
  END TX_BIAS_I[1]
  PIN RX_GAIN_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8075 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.036 LAYER C2 ;
      ANTENNAMAXAREACAR 346.412778 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 87.71 80 87.87 ;
    END
  END RX_GAIN_I[3]
  PIN TX_BIAS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 153.23 80 153.39 ;
    END
  END TX_BIAS_I[3]
  PIN DI_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2128 LAYER C2 ;
    ANTENNADIFFAREA 0.16192 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 129.83 80 129.99 ;
    END
  END DI_O
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2128 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C2 ;
      ANTENNAMAXAREACAR 30.536607 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 130.87 80 131.03 ;
    END
  END DO_I
  PIN EI_DETECT_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2128 LAYER C2 ;
    ANTENNADIFFAREA 0.081 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 49.23 80 49.39 ;
    END
  END EI_DETECT_O
  PIN RX_CTLE_RES_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8075 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0198 LAYER C2 ;
      ANTENNAMAXAREACAR 470.405051 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 92.13 80 92.29 ;
    END
  END RX_CTLE_RES_I[4]
  PIN RTERM_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 28.891274 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 175.07 80 175.23 ;
    END
  END RTERM_EN_I
  PIN RTERM_TRIM_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 175.59 80 175.75 ;
    END
  END RTERM_TRIM_I[0]
  PIN RTERM_TRIM_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 176.11 80 176.27 ;
    END
  END RTERM_TRIM_I[1]
  PIN RTERM_TRIM_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 176.63 80 176.79 ;
    END
  END RTERM_TRIM_I[2]
  PIN RTERM_TRIM_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 177.15 80 177.31 ;
    END
  END RTERM_TRIM_I[3]
  PIN RX_POL_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0224 LAYER C2 ;
      ANTENNAMAXAREACAR 56.869643 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 128.27 80 128.43 ;
    END
  END RX_POL_I
  PIN TX_FFE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23216 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02128 LAYER C2 ;
      ANTENNAMAXAREACAR 26.403195 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 129.31 80 129.47 ;
    END
  END TX_FFE_I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 64.05 0 67.65 180 ;
    END
    PORT
      LAYER JA ;
        RECT 68.75 0 72.35 180 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 166.05 80 169.05 ;
      LAYER OI ;
        RECT 78.15 166.05 80 169.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 161.35 80 164.35 ;
      LAYER OI ;
        RECT 78.15 161.35 80 164.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 147.25 80 150.25 ;
      LAYER OI ;
        RECT 78.15 147.25 80 150.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 142.55 80 145.55 ;
      LAYER OI ;
        RECT 78.15 142.55 80 145.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 128.45 80 131.45 ;
      LAYER OI ;
        RECT 78.15 128.45 80 131.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 123.75 80 126.75 ;
      LAYER OI ;
        RECT 78.15 123.75 80 126.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 109.65 80 112.65 ;
      LAYER OI ;
        RECT 78.15 109.65 80 112.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 104.95 80 107.95 ;
      LAYER OI ;
        RECT 78.15 104.95 80 107.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 90.85 80 93.85 ;
      LAYER OI ;
        RECT 78.15 90.85 80 93.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 86.15 80 89.15 ;
      LAYER OI ;
        RECT 78.15 86.15 80 89.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 72.05 80 75.05 ;
      LAYER OI ;
        RECT 78.15 72.05 80 75.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 67.35 80 70.35 ;
      LAYER OI ;
        RECT 78.15 67.35 80 70.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 53.25 80 56.25 ;
      LAYER OI ;
        RECT 78.15 53.25 80 56.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 48.55 80 51.55 ;
      LAYER OI ;
        RECT 78.15 48.55 80 51.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 34.45 80 37.45 ;
      LAYER OI ;
        RECT 78.15 34.45 80 37.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 29.75 80 32.75 ;
      LAYER OI ;
        RECT 78.15 29.75 80 32.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 15.65 80 18.65 ;
      LAYER OI ;
        RECT 78.15 15.65 80 18.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 10.95 80 13.95 ;
      LAYER OI ;
        RECT 78.15 10.95 80 13.95 ;
    END
  END VDD
  PIN TX_EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34096 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 28.164002 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 151.15 80 151.31 ;
    END
  END TX_EN_I
  OBS
    LAYER CA ;
      RECT 0 0 80 180 ;
    LAYER M1 ;
      RECT 0 0 80 180 ;
    LAYER V1 ;
      RECT 0 0 80 180 ;
    LAYER M2 ;
      RECT 0 0 80 180 ;
    LAYER A1 ;
      RECT 0 0 80 180 ;
    LAYER C2 ;
      RECT 0 0 80 180 ;
    LAYER CB ;
      RECT 0 0 80 180 ;
    LAYER YS ;
      RECT 0 0 80 180 ;
    LAYER OI ;
      RECT 0 0 80 180 ;
    LAYER JQ ;
      RECT 0 0 80 180 ;
    LAYER JA ;
      RECT 0 0 80 180 ;
    LAYER AY ;
      RECT 0 0 80 180 ;
    LAYER C1 ;
      RECT 0 0 80 180 ;
    LAYER C5 ;
      RECT 0 0 80 180 ;
    LAYER C4 ;
      RECT 0 0 80 180 ;
    LAYER C3 ;
      RECT 0 0 80 180 ;
    LAYER A4 ;
      RECT 0 0 80 180 ;
    LAYER A3 ;
      RECT 0 0 80 180 ;
    LAYER A2 ;
      RECT 0 0 80 180 ;
  END
END RIIO_EG1D80V_HPLVDS_TX_SLVT28_H

MACRO RIIO_EG1D80V_RTERMCAL_HVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_HVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER JA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER JA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER JA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER JA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER JA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER JA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER JA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.46 80 40.6 ;
    END
  END VSSQ
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER JA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER JA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER JA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER JA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.8325 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER JA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 48.28176 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 9.405088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 15.42564 LAYER YS ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.663328 LAYER A2 ;
    ANTENNADIFFAREA 152.2484 LAYER C4 ;
    ANTENNADIFFAREA 152.2484 LAYER C3 ;
    ANTENNADIFFAREA 152.2484 LAYER C5 ;
    ANTENNADIFFAREA 152.2484 LAYER JA ;
    ANTENNADIFFAREA 152.2484 LAYER OI ;
    ANTENNADIFFAREA 152.2484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER JA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 98.217391 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.74 80 47.88 ;
    END
  END MODE_I[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 52.609456 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.22 80 47.36 ;
    END
  END MODE_I[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.7 80 46.84 ;
    END
  END RESULT_O[0]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.18 80 46.32 ;
    END
  END RESULT_O[1]
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.02 80 55.16 ;
    END
  END D_IOSG_I[10]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.811972 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.54 80 55.68 ;
    END
  END D_IOSG_I[11]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.82975 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.06 80 56.2 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C2 ;
      ANTENNAMAXAREACAR 14.865466 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.58 80 56.72 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C2 ;
      ANTENNAMAXAREACAR 14.455976 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.1 80 57.24 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C2 ;
      ANTENNAMAXAREACAR 13.688986 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.62 80 57.76 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.665245 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.34 80 50.48 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.666814 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.86 80 51 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.38 80 51.52 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.9 80 52.04 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.42 80 52.56 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.94 80 53.08 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.46 80 53.6 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.98 80 54.12 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 54.5 80 54.64 ;
    END
  END D_IOSG_I[9]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.629464 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.82 80 49.96 ;
    END
  END D_LVDS_I[0]
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.950893 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.3 80 49.44 ;
    END
  END D_LVDS_I[1]
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.98 80 41.12 ;
    END
  END VDDQ
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.236607 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.78 80 48.92 ;
    END
  END D_LVDS_I[2]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.558036 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.26 80 48.4 ;
    END
  END D_LVDS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_RTERMCAL_HVT28_H

MACRO RIIO_EG1D80V_RTERMCAL_LLHVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_LLHVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER JA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER JA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER JA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER JA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER JA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER JA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER JA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.46 80 40.6 ;
    END
  END VSSQ
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER JA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER JA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER JA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER JA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.8325 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER JA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 48.28176 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 9.405088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 15.42564 LAYER YS ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.663328 LAYER A2 ;
    ANTENNADIFFAREA 152.2484 LAYER C4 ;
    ANTENNADIFFAREA 152.2484 LAYER C3 ;
    ANTENNADIFFAREA 152.2484 LAYER C5 ;
    ANTENNADIFFAREA 152.2484 LAYER JA ;
    ANTENNADIFFAREA 152.2484 LAYER OI ;
    ANTENNADIFFAREA 152.2484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER JA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0184 LAYER C2 ;
      ANTENNAMAXAREACAR 138.063043 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.74 80 47.88 ;
    END
  END MODE_I[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.044 LAYER C2 ;
      ANTENNAMAXAREACAR 72.110568 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.22 80 47.36 ;
    END
  END MODE_I[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.03864 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.7 80 46.84 ;
    END
  END RESULT_O[0]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.03864 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.18 80 46.32 ;
    END
  END RESULT_O[1]
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.02 80 55.16 ;
    END
  END D_IOSG_I[10]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.811972 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.54 80 55.68 ;
    END
  END D_IOSG_I[11]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.82975 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.06 80 56.2 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C2 ;
      ANTENNAMAXAREACAR 14.865466 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.58 80 56.72 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C2 ;
      ANTENNAMAXAREACAR 14.455976 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.1 80 57.24 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C2 ;
      ANTENNAMAXAREACAR 13.688986 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.62 80 57.76 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.665245 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.34 80 50.48 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.666814 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.86 80 51 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.38 80 51.52 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.9 80 52.04 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.42 80 52.56 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.94 80 53.08 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.46 80 53.6 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.98 80 54.12 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 54.5 80 54.64 ;
    END
  END D_IOSG_I[9]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C2 ;
      ANTENNAMAXAREACAR 399.80625 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.82 80 49.96 ;
    END
  END D_LVDS_I[0]
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C2 ;
      ANTENNAMAXAREACAR 399.15625 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.3 80 49.44 ;
    END
  END D_LVDS_I[1]
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.98 80 41.12 ;
    END
  END VDDQ
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C2 ;
      ANTENNAMAXAREACAR 399.15625 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.78 80 48.92 ;
    END
  END D_LVDS_I[2]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0064 LAYER C2 ;
      ANTENNAMAXAREACAR 399.15625 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.26 80 48.4 ;
    END
  END D_LVDS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_RTERMCAL_LLHVT28_H

MACRO RIIO_EG1D80V_RTERMCAL_LVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_LVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER JA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER JA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER JA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER JA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER JA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER JA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER JA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.46 80 40.6 ;
    END
  END VSSQ
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER JA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER JA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER JA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER JA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.8325 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER JA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 48.28176 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 9.405088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 15.42564 LAYER YS ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.663328 LAYER A2 ;
    ANTENNADIFFAREA 152.2484 LAYER C4 ;
    ANTENNADIFFAREA 152.2484 LAYER C3 ;
    ANTENNADIFFAREA 152.2484 LAYER C5 ;
    ANTENNADIFFAREA 152.2484 LAYER JA ;
    ANTENNADIFFAREA 152.2484 LAYER OI ;
    ANTENNADIFFAREA 152.2484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER JA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 98.217391 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.74 80 47.88 ;
    END
  END MODE_I[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 52.609456 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.22 80 47.36 ;
    END
  END MODE_I[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.7 80 46.84 ;
    END
  END RESULT_O[0]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.18 80 46.32 ;
    END
  END RESULT_O[1]
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.02 80 55.16 ;
    END
  END D_IOSG_I[10]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.811972 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.54 80 55.68 ;
    END
  END D_IOSG_I[11]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.82975 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.06 80 56.2 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C2 ;
      ANTENNAMAXAREACAR 14.865466 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.58 80 56.72 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C2 ;
      ANTENNAMAXAREACAR 14.455976 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.1 80 57.24 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C2 ;
      ANTENNAMAXAREACAR 13.688986 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.62 80 57.76 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.665245 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.34 80 50.48 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.666814 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.86 80 51 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.38 80 51.52 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.9 80 52.04 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.42 80 52.56 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.94 80 53.08 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.46 80 53.6 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.98 80 54.12 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 54.5 80 54.64 ;
    END
  END D_IOSG_I[9]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.629464 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.82 80 49.96 ;
    END
  END D_LVDS_I[0]
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.950893 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.3 80 49.44 ;
    END
  END D_LVDS_I[1]
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.98 80 41.12 ;
    END
  END VDDQ
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.236607 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.78 80 48.92 ;
    END
  END D_LVDS_I[2]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.558036 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.26 80 48.4 ;
    END
  END D_LVDS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_RTERMCAL_LVT28_H

MACRO RIIO_EG1D80V_RTERMCAL_RVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER JA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER JA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER JA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER JA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER JA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER JA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER JA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.46 80 40.6 ;
    END
  END VSSQ
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER JA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER JA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER JA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER JA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.8325 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER JA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 48.28176 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 9.405088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 15.42564 LAYER YS ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.663328 LAYER A2 ;
    ANTENNADIFFAREA 152.2484 LAYER C4 ;
    ANTENNADIFFAREA 152.2484 LAYER C3 ;
    ANTENNADIFFAREA 152.2484 LAYER C5 ;
    ANTENNADIFFAREA 152.2484 LAYER JA ;
    ANTENNADIFFAREA 152.2484 LAYER OI ;
    ANTENNADIFFAREA 152.2484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER JA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 98.217391 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.74 80 47.88 ;
    END
  END MODE_I[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 52.609456 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.22 80 47.36 ;
    END
  END MODE_I[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.7 80 46.84 ;
    END
  END RESULT_O[0]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.18 80 46.32 ;
    END
  END RESULT_O[1]
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.02 80 55.16 ;
    END
  END D_IOSG_I[10]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.811972 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.54 80 55.68 ;
    END
  END D_IOSG_I[11]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.82975 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.06 80 56.2 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C2 ;
      ANTENNAMAXAREACAR 14.865466 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.58 80 56.72 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C2 ;
      ANTENNAMAXAREACAR 14.455976 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.1 80 57.24 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C2 ;
      ANTENNAMAXAREACAR 13.688986 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.62 80 57.76 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.665245 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.34 80 50.48 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.666814 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.86 80 51 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.38 80 51.52 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.9 80 52.04 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.42 80 52.56 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.94 80 53.08 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.46 80 53.6 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.98 80 54.12 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 54.5 80 54.64 ;
    END
  END D_IOSG_I[9]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.629464 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.82 80 49.96 ;
    END
  END D_LVDS_I[0]
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.950893 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.3 80 49.44 ;
    END
  END D_LVDS_I[1]
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.98 80 41.12 ;
    END
  END VDDQ
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.236607 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.78 80 48.92 ;
    END
  END D_LVDS_I[2]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.558036 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.26 80 48.4 ;
    END
  END D_LVDS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_RTERMCAL_RVT28_H

MACRO RIIO_EG1D80V_RTERMCAL_SLVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RTERMCAL_SLVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER JA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER JA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER JA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER JA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER JA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER JA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER JA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER JA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER JA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER JA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER JA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.46 80 40.6 ;
    END
  END VSSQ
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER JA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER JA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER JA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER JA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER JA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.8325 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER JA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 48.28176 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 9.405088 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 15.42564 LAYER YS ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.663328 LAYER A2 ;
    ANTENNADIFFAREA 152.2484 LAYER C4 ;
    ANTENNADIFFAREA 152.2484 LAYER C3 ;
    ANTENNADIFFAREA 152.2484 LAYER C5 ;
    ANTENNADIFFAREA 152.2484 LAYER JA ;
    ANTENNADIFFAREA 152.2484 LAYER OI ;
    ANTENNADIFFAREA 152.2484 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER JA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN MODE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 98.217391 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.74 80 47.88 ;
    END
  END MODE_I[0]
  PIN MODE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0616 LAYER C2 ;
      ANTENNAMAXAREACAR 52.609456 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 47.22 80 47.36 ;
    END
  END MODE_I[1]
  PIN RESULT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.7 80 46.84 ;
    END
  END RESULT_O[0]
  PIN RESULT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 46.18 80 46.32 ;
    END
  END RESULT_O[1]
  PIN D_IOSG_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.02 80 55.16 ;
    END
  END D_IOSG_I[10]
  PIN D_IOSG_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.811972 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 55.54 80 55.68 ;
    END
  END D_IOSG_I[11]
  PIN D_IOSG_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER C2 ;
      ANTENNAMAXAREACAR 16.82975 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.06 80 56.2 ;
    END
  END D_IOSG_I[12]
  PIN D_IOSG_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.408 LAYER C2 ;
      ANTENNAMAXAREACAR 14.865466 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 56.58 80 56.72 ;
    END
  END D_IOSG_I[13]
  PIN D_IOSG_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.42 LAYER C2 ;
      ANTENNAMAXAREACAR 14.455976 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.1 80 57.24 ;
    END
  END D_IOSG_I[14]
  PIN D_IOSG_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.444 LAYER C2 ;
      ANTENNAMAXAREACAR 13.688986 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 57.62 80 57.76 ;
    END
  END D_IOSG_I[15]
  PIN D_IOSG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.665245 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.34 80 50.48 ;
    END
  END D_IOSG_I[1]
  PIN D_IOSG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.204 LAYER C2 ;
      ANTENNAMAXAREACAR 29.666814 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 50.86 80 51 ;
    END
  END D_IOSG_I[2]
  PIN D_IOSG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.38 80 51.52 ;
    END
  END D_IOSG_I[3]
  PIN D_IOSG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER C2 ;
      ANTENNAMAXAREACAR 28.009769 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 51.9 80 52.04 ;
    END
  END D_IOSG_I[4]
  PIN D_IOSG_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.42 80 52.56 ;
    END
  END D_IOSG_I[5]
  PIN D_IOSG_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER C2 ;
      ANTENNAMAXAREACAR 25.208792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 52.94 80 53.08 ;
    END
  END D_IOSG_I[6]
  PIN D_IOSG_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.46 80 53.6 ;
    END
  END D_IOSG_I[7]
  PIN D_IOSG_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER C2 ;
      ANTENNAMAXAREACAR 21.920688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 53.98 80 54.12 ;
    END
  END D_IOSG_I[8]
  PIN D_IOSG_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.336 LAYER C2 ;
      ANTENNAMAXAREACAR 18.00628 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 54.5 80 54.64 ;
    END
  END D_IOSG_I[9]
  PIN D_LVDS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.629464 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.82 80 49.96 ;
    END
  END D_LVDS_I[0]
  PIN D_LVDS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.950893 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 49.3 80 49.44 ;
    END
  END D_LVDS_I[1]
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 79.86 40.98 80 41.12 ;
    END
  END VDDQ
  PIN D_LVDS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.236607 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.78 80 48.92 ;
    END
  END D_LVDS_I[2]
  PIN D_LVDS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00896 LAYER C2 ;
      ANTENNAMAXAREACAR 286.558036 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.86 48.26 80 48.4 ;
    END
  END D_LVDS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_RTERMCAL_SLVT28_H

END LIBRARY
