VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RIIO_EG1D80V_CORNER_45
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CORNER_45 0 0 ;
  SIZE 80 BY 80 ;
  SYMMETRY X Y ;
  SITE corner_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 75.44 61.2 80 66 ;
        RECT 70.646 65.971 77.43 66.006 ;
        RECT 68.668 67.949 75.44 67.995 ;
        RECT 68.714 67.903 75.486 67.967 ;
        RECT 75.43 61.205 75.44 67.995 ;
        RECT 68.76 67.857 75.532 67.921 ;
        RECT 75.384 61.233 75.43 68.023 ;
        RECT 68.622 67.995 75.384 68.069 ;
        RECT 68.806 67.811 75.578 67.875 ;
        RECT 75.338 61.279 75.384 68.069 ;
        RECT 68.576 68.041 75.338 68.115 ;
        RECT 68.852 67.765 75.624 67.829 ;
        RECT 75.292 61.325 75.338 68.115 ;
        RECT 68.53 68.087 75.292 68.161 ;
        RECT 68.898 67.719 75.67 67.783 ;
        RECT 75.246 61.371 75.292 68.161 ;
        RECT 68.484 68.133 75.246 68.207 ;
        RECT 68.944 67.673 75.716 67.737 ;
        RECT 75.2 61.417 75.246 68.207 ;
        RECT 68.438 68.179 75.2 68.253 ;
        RECT 68.99 67.627 75.762 67.691 ;
        RECT 75.154 61.463 75.2 68.253 ;
        RECT 68.392 68.225 75.154 68.299 ;
        RECT 69.036 67.581 75.808 67.645 ;
        RECT 75.108 61.509 75.154 68.299 ;
        RECT 68.346 68.271 75.108 68.345 ;
        RECT 69.082 67.535 75.854 67.599 ;
        RECT 75.062 61.555 75.108 68.345 ;
        RECT 68.3 68.317 75.062 68.391 ;
        RECT 69.128 67.489 75.9 67.553 ;
        RECT 75.016 61.601 75.062 68.391 ;
        RECT 68.254 68.363 75.016 68.437 ;
        RECT 69.174 67.443 75.946 67.507 ;
        RECT 74.97 61.647 75.016 68.437 ;
        RECT 68.208 68.409 74.97 68.483 ;
        RECT 69.22 67.397 75.992 67.461 ;
        RECT 74.924 61.693 74.97 68.483 ;
        RECT 68.162 68.455 74.924 68.529 ;
        RECT 69.266 67.351 76.038 67.415 ;
        RECT 74.878 61.739 74.924 68.529 ;
        RECT 68.116 68.501 74.878 68.575 ;
        RECT 69.312 67.305 76.084 67.369 ;
        RECT 74.832 61.785 74.878 68.575 ;
        RECT 68.07 68.547 74.832 68.621 ;
        RECT 69.358 67.259 76.13 67.323 ;
        RECT 74.786 61.831 74.832 68.621 ;
        RECT 68.024 68.593 74.786 68.667 ;
        RECT 69.404 67.213 76.176 67.277 ;
        RECT 74.74 61.877 74.786 68.667 ;
        RECT 67.978 68.639 74.74 68.713 ;
        RECT 69.45 67.167 76.222 67.231 ;
        RECT 74.694 61.923 74.74 68.713 ;
        RECT 67.932 68.685 74.694 68.759 ;
        RECT 69.496 67.121 76.268 67.185 ;
        RECT 74.648 61.969 74.694 68.759 ;
        RECT 67.886 68.731 74.648 68.805 ;
        RECT 69.542 67.075 76.314 67.139 ;
        RECT 74.602 62.015 74.648 68.805 ;
        RECT 67.84 68.777 74.602 68.851 ;
        RECT 69.588 67.029 76.36 67.093 ;
        RECT 74.556 62.061 74.602 68.851 ;
        RECT 67.794 68.823 74.556 68.897 ;
        RECT 69.634 66.983 76.406 67.047 ;
        RECT 74.51 62.107 74.556 68.897 ;
        RECT 67.748 68.869 74.51 68.943 ;
        RECT 69.68 66.937 76.452 67.001 ;
        RECT 74.464 62.153 74.51 68.943 ;
        RECT 67.702 68.915 74.464 68.989 ;
        RECT 69.726 66.891 76.498 66.955 ;
        RECT 74.418 62.199 74.464 68.989 ;
        RECT 67.656 68.961 74.418 69.035 ;
        RECT 69.772 66.845 76.544 66.909 ;
        RECT 74.372 62.245 74.418 69.035 ;
        RECT 67.61 69.007 74.372 69.081 ;
        RECT 69.818 66.799 76.59 66.863 ;
        RECT 74.326 62.291 74.372 69.081 ;
        RECT 67.564 69.053 74.326 69.127 ;
        RECT 69.864 66.753 76.636 66.817 ;
        RECT 74.28 62.337 74.326 69.127 ;
        RECT 67.518 69.099 74.28 69.173 ;
        RECT 69.91 66.707 76.682 66.771 ;
        RECT 74.234 62.383 74.28 69.173 ;
        RECT 67.472 69.145 74.234 69.219 ;
        RECT 69.956 66.661 76.728 66.725 ;
        RECT 74.188 62.429 74.234 69.219 ;
        RECT 67.426 69.191 74.188 69.265 ;
        RECT 70.002 66.615 76.774 66.679 ;
        RECT 74.142 62.475 74.188 69.265 ;
        RECT 67.38 69.237 74.142 69.311 ;
        RECT 70.048 66.569 76.82 66.633 ;
        RECT 74.096 62.521 74.142 69.311 ;
        RECT 67.334 69.283 74.096 69.357 ;
        RECT 70.094 66.523 76.866 66.587 ;
        RECT 74.05 62.567 74.096 69.357 ;
        RECT 67.288 69.329 74.05 69.403 ;
        RECT 70.14 66.477 76.912 66.541 ;
        RECT 74.004 62.613 74.05 69.403 ;
        RECT 67.242 69.375 74.004 69.449 ;
        RECT 70.186 66.431 76.958 66.495 ;
        RECT 73.958 62.659 74.004 69.449 ;
        RECT 67.196 69.421 73.958 69.495 ;
        RECT 70.232 66.385 77.004 66.449 ;
        RECT 73.912 62.705 73.958 69.495 ;
        RECT 67.15 69.467 73.912 69.541 ;
        RECT 70.278 66.339 77.05 66.403 ;
        RECT 73.866 62.751 73.912 69.541 ;
        RECT 67.104 69.513 73.866 69.587 ;
        RECT 70.324 66.293 77.096 66.357 ;
        RECT 73.82 62.797 73.866 69.587 ;
        RECT 67.058 69.559 73.82 69.633 ;
        RECT 70.37 66.247 77.142 66.311 ;
        RECT 73.774 62.843 73.82 69.633 ;
        RECT 67.012 69.605 73.774 69.679 ;
        RECT 70.416 66.201 77.188 66.265 ;
        RECT 73.728 62.889 73.774 69.679 ;
        RECT 66.966 69.651 73.728 69.725 ;
        RECT 70.462 66.155 77.234 66.219 ;
        RECT 73.682 62.935 73.728 69.725 ;
        RECT 66.92 69.697 73.682 69.771 ;
        RECT 70.508 66.109 77.28 66.173 ;
        RECT 73.636 62.981 73.682 69.771 ;
        RECT 66.874 69.743 73.636 69.817 ;
        RECT 70.554 66.063 77.326 66.127 ;
        RECT 73.59 63.027 73.636 69.817 ;
        RECT 66.828 69.789 73.59 69.863 ;
        RECT 70.6 66.017 77.372 66.081 ;
        RECT 73.544 63.073 73.59 69.863 ;
        RECT 66.782 69.835 73.544 69.909 ;
        RECT 70.646 65.971 77.418 66.035 ;
        RECT 73.498 63.119 73.544 69.909 ;
        RECT 66.736 69.881 73.498 69.955 ;
        RECT 70.692 65.925 80 66 ;
        RECT 73.452 63.165 73.498 69.955 ;
        RECT 66.69 69.927 73.452 70.001 ;
        RECT 70.738 65.879 80 66 ;
        RECT 73.406 63.211 73.452 70.001 ;
        RECT 66.644 69.973 73.406 70.047 ;
        RECT 70.784 65.833 80 66 ;
        RECT 73.36 63.257 73.406 70.047 ;
        RECT 66.598 70.019 73.36 70.093 ;
        RECT 70.83 65.787 80 66 ;
        RECT 73.314 63.303 73.36 70.093 ;
        RECT 66.552 70.065 73.314 70.139 ;
        RECT 70.876 65.741 80 66 ;
        RECT 73.268 63.349 73.314 70.139 ;
        RECT 66.506 70.111 73.268 70.185 ;
        RECT 70.922 65.695 80 66 ;
        RECT 73.222 63.395 73.268 70.185 ;
        RECT 66.46 70.157 73.222 70.231 ;
        RECT 70.968 65.649 80 66 ;
        RECT 73.176 63.441 73.222 70.231 ;
        RECT 66.414 70.203 73.176 70.277 ;
        RECT 71.014 65.603 80 66 ;
        RECT 73.13 63.487 73.176 70.277 ;
        RECT 66.368 70.249 73.13 70.323 ;
        RECT 71.06 65.557 80 66 ;
        RECT 73.084 63.533 73.13 70.323 ;
        RECT 66.322 70.295 73.084 70.369 ;
        RECT 71.106 65.511 80 66 ;
        RECT 73.038 63.579 73.084 70.369 ;
        RECT 66.276 70.341 73.038 70.415 ;
        RECT 71.152 65.465 80 66 ;
        RECT 72.992 63.625 73.038 70.415 ;
        RECT 66.23 70.387 72.992 70.461 ;
        RECT 71.198 65.419 80 66 ;
        RECT 72.946 63.671 72.992 70.461 ;
        RECT 66.184 70.433 72.946 70.507 ;
        RECT 71.244 65.373 80 66 ;
        RECT 72.9 63.717 72.946 70.507 ;
        RECT 66.138 70.479 72.9 70.553 ;
        RECT 71.29 65.327 80 66 ;
        RECT 72.854 63.763 72.9 70.553 ;
        RECT 66.092 70.525 72.854 70.599 ;
        RECT 71.336 65.281 80 66 ;
        RECT 72.808 63.809 72.854 70.599 ;
        RECT 66.046 70.571 72.808 70.645 ;
        RECT 71.382 65.235 80 66 ;
        RECT 72.762 63.855 72.808 70.645 ;
        RECT 65.984 70.648 72.762 70.691 ;
        RECT 66 70.617 72.762 70.691 ;
        RECT 71.428 65.189 80 66 ;
        RECT 72.716 63.901 72.762 70.691 ;
        RECT 65.938 70.679 72.716 70.737 ;
        RECT 71.474 65.143 80 66 ;
        RECT 72.67 63.947 72.716 70.737 ;
        RECT 65.892 70.725 72.67 70.783 ;
        RECT 71.52 65.097 80 66 ;
        RECT 72.624 63.993 72.67 70.783 ;
        RECT 65.846 70.771 72.624 70.829 ;
        RECT 71.566 65.051 80 66 ;
        RECT 72.578 64.039 72.624 70.829 ;
        RECT 65.8 70.817 72.578 70.875 ;
        RECT 71.612 65.005 80 66 ;
        RECT 72.532 64.085 72.578 70.875 ;
        RECT 65.754 70.863 72.532 70.921 ;
        RECT 71.658 64.959 80 66 ;
        RECT 72.486 64.131 72.532 70.921 ;
        RECT 65.708 70.909 72.486 70.967 ;
        RECT 71.704 64.913 80 66 ;
        RECT 72.44 64.177 72.486 70.967 ;
        RECT 65.662 70.955 72.44 71.013 ;
        RECT 71.75 64.867 80 66 ;
        RECT 72.394 64.223 72.44 71.013 ;
        RECT 65.616 71.001 72.394 71.059 ;
        RECT 71.796 64.821 80 66 ;
        RECT 72.348 64.269 72.394 71.059 ;
        RECT 65.57 71.047 72.348 71.105 ;
        RECT 71.842 64.775 80 66 ;
        RECT 72.302 64.315 72.348 71.105 ;
        RECT 65.524 71.093 72.302 71.151 ;
        RECT 71.888 64.729 80 66 ;
        RECT 72.256 64.361 72.302 71.151 ;
        RECT 65.478 71.139 72.256 71.197 ;
        RECT 71.934 64.683 80 66 ;
        RECT 72.21 64.407 72.256 71.197 ;
        RECT 65.432 71.185 72.21 71.243 ;
        RECT 71.98 64.637 80 66 ;
        RECT 72.164 64.453 72.21 71.243 ;
        RECT 65.386 71.231 72.164 71.289 ;
        RECT 72.026 64.591 80 66 ;
        RECT 72.118 64.499 72.164 71.289 ;
        RECT 65.34 71.277 72.118 71.335 ;
        RECT 72.072 64.545 80 66 ;
        RECT 65.294 71.323 72.072 71.381 ;
        RECT 65.248 71.369 72.026 71.427 ;
        RECT 65.202 71.415 71.98 71.473 ;
        RECT 65.156 71.461 71.934 71.519 ;
        RECT 65.11 71.507 71.888 71.565 ;
        RECT 65.064 71.553 71.842 71.611 ;
        RECT 65.018 71.599 71.796 71.657 ;
        RECT 64.972 71.645 71.75 71.703 ;
        RECT 64.926 71.691 71.704 71.749 ;
        RECT 64.88 71.737 71.658 71.795 ;
        RECT 64.834 71.783 71.612 71.841 ;
        RECT 64.788 71.829 71.566 71.887 ;
        RECT 64.742 71.875 71.52 71.933 ;
        RECT 64.696 71.921 71.474 71.979 ;
        RECT 64.65 71.967 71.428 72.025 ;
        RECT 64.604 72.013 71.382 72.071 ;
        RECT 64.558 72.059 71.336 72.117 ;
        RECT 64.512 72.105 71.29 72.163 ;
        RECT 64.466 72.151 71.244 72.209 ;
        RECT 64.42 72.197 71.198 72.255 ;
        RECT 64.374 72.243 71.152 72.301 ;
        RECT 64.328 72.289 71.106 72.347 ;
        RECT 64.282 72.335 71.06 72.393 ;
        RECT 64.236 72.381 71.014 72.439 ;
        RECT 64.19 72.427 70.968 72.485 ;
        RECT 64.144 72.473 70.922 72.531 ;
        RECT 64.098 72.519 70.876 72.577 ;
        RECT 64.052 72.565 70.83 72.623 ;
        RECT 64.006 72.611 70.784 72.669 ;
        RECT 63.96 72.657 70.738 72.715 ;
        RECT 63.914 72.703 70.692 72.761 ;
        RECT 63.868 72.749 70.646 72.807 ;
        RECT 63.822 72.795 70.6 72.853 ;
        RECT 63.776 72.841 70.554 72.899 ;
        RECT 63.73 72.887 70.508 72.945 ;
        RECT 63.684 72.933 70.462 72.991 ;
        RECT 63.638 72.979 70.416 73.037 ;
        RECT 63.592 73.025 70.37 73.083 ;
        RECT 63.546 73.071 70.324 73.129 ;
        RECT 63.5 73.117 70.278 73.175 ;
        RECT 63.454 73.163 70.232 73.221 ;
        RECT 63.408 73.209 70.186 73.267 ;
        RECT 63.362 73.255 70.14 73.313 ;
        RECT 63.316 73.301 70.094 73.359 ;
        RECT 63.27 73.347 70.048 73.405 ;
        RECT 63.224 73.393 70.002 73.451 ;
        RECT 63.178 73.439 69.956 73.497 ;
        RECT 63.132 73.485 69.91 73.543 ;
        RECT 63.086 73.531 69.864 73.589 ;
        RECT 63.04 73.577 69.818 73.635 ;
        RECT 62.994 73.623 69.772 73.681 ;
        RECT 62.948 73.669 69.726 73.727 ;
        RECT 62.902 73.715 69.68 73.773 ;
        RECT 62.856 73.761 69.634 73.819 ;
        RECT 62.81 73.807 69.588 73.865 ;
        RECT 62.764 73.853 69.542 73.911 ;
        RECT 62.718 73.899 69.496 73.957 ;
        RECT 62.672 73.945 69.45 74.003 ;
        RECT 62.626 73.991 69.404 74.049 ;
        RECT 62.58 74.037 69.358 74.095 ;
        RECT 62.534 74.083 69.312 74.141 ;
        RECT 62.488 74.129 69.266 74.187 ;
        RECT 62.442 74.175 69.22 74.233 ;
        RECT 62.396 74.221 69.174 74.279 ;
        RECT 62.35 74.267 69.128 74.325 ;
        RECT 62.304 74.313 69.082 74.371 ;
        RECT 62.258 74.359 69.036 74.417 ;
        RECT 62.212 74.405 68.99 74.463 ;
        RECT 62.166 74.451 68.944 74.509 ;
        RECT 62.12 74.497 68.898 74.555 ;
        RECT 62.074 74.543 68.852 74.601 ;
        RECT 62.028 74.589 68.806 74.647 ;
        RECT 61.982 74.635 68.76 74.693 ;
        RECT 61.936 74.681 68.714 74.739 ;
        RECT 61.89 74.727 68.668 74.785 ;
        RECT 61.844 74.773 68.622 74.831 ;
        RECT 61.798 74.819 68.576 74.877 ;
        RECT 61.752 74.865 68.53 74.923 ;
        RECT 61.706 74.911 68.484 74.969 ;
        RECT 61.66 74.957 68.438 75.015 ;
        RECT 61.614 75.003 68.392 75.061 ;
        RECT 61.568 75.049 68.346 75.107 ;
        RECT 61.522 75.095 68.3 75.153 ;
        RECT 61.476 75.141 68.254 75.199 ;
        RECT 61.43 75.187 68.208 75.245 ;
        RECT 61.384 75.233 68.162 75.291 ;
        RECT 61.338 75.279 68.116 75.337 ;
        RECT 61.292 75.325 68.07 75.383 ;
        RECT 61.246 75.371 68.024 75.429 ;
        RECT 61.2 75.417 67.978 75.475 ;
        RECT 61.2 75.417 67.932 75.521 ;
        RECT 61.2 75.417 67.886 75.567 ;
        RECT 61.2 75.417 67.84 75.613 ;
        RECT 61.2 75.417 67.794 75.659 ;
        RECT 61.2 75.417 67.748 75.705 ;
        RECT 61.2 75.417 67.702 75.751 ;
        RECT 61.2 75.417 67.656 75.797 ;
        RECT 61.2 75.417 67.61 75.843 ;
        RECT 61.2 75.417 67.564 75.889 ;
        RECT 61.2 75.417 67.518 75.935 ;
        RECT 61.2 75.417 67.472 75.981 ;
        RECT 61.2 75.417 67.426 76.027 ;
        RECT 61.2 75.417 67.38 76.073 ;
        RECT 61.2 75.417 67.334 76.119 ;
        RECT 61.2 75.417 67.288 76.165 ;
        RECT 61.2 75.417 67.242 76.211 ;
        RECT 61.2 75.417 67.196 76.257 ;
        RECT 61.2 75.417 67.15 76.303 ;
        RECT 61.2 75.417 67.104 76.349 ;
        RECT 61.2 75.417 67.058 76.395 ;
        RECT 61.2 75.417 67.012 76.441 ;
        RECT 61.2 75.417 66.966 76.487 ;
        RECT 61.2 75.417 66.92 76.533 ;
        RECT 61.2 75.417 66.874 76.579 ;
        RECT 61.2 75.417 66.828 76.625 ;
        RECT 61.2 75.417 66.782 76.671 ;
        RECT 61.2 75.417 66.736 76.717 ;
        RECT 61.2 75.417 66.69 76.763 ;
        RECT 61.2 75.417 66.644 76.809 ;
        RECT 61.2 75.417 66.598 76.855 ;
        RECT 61.2 75.417 66.552 76.901 ;
        RECT 61.2 75.417 66.506 76.947 ;
        RECT 61.2 75.417 66.46 76.993 ;
        RECT 61.2 75.417 66.414 77.039 ;
        RECT 61.2 75.417 66.368 77.085 ;
        RECT 61.2 75.417 66.322 77.131 ;
        RECT 61.2 75.417 66.276 77.177 ;
        RECT 61.2 75.417 66.23 77.223 ;
        RECT 61.2 75.417 66.184 77.269 ;
        RECT 61.2 75.417 66.138 77.315 ;
        RECT 61.2 75.417 66.092 77.361 ;
        RECT 61.2 75.417 66.046 77.407 ;
        RECT 61.2 75.417 66 80 ;
    END
    PORT
      LAYER QB ;
        RECT 72.87 55 80 59.8 ;
        RECT 68.08 59.767 74.86 59.806 ;
        RECT 66.102 61.745 72.87 61.793 ;
        RECT 66.148 61.699 72.916 61.767 ;
        RECT 72.864 55.003 72.87 61.793 ;
        RECT 66.194 61.653 72.962 61.721 ;
        RECT 72.818 55.029 72.864 61.819 ;
        RECT 66.056 61.791 72.818 61.865 ;
        RECT 66.24 61.607 73.008 61.675 ;
        RECT 72.772 55.075 72.818 61.865 ;
        RECT 66.01 61.837 72.772 61.911 ;
        RECT 66.286 61.561 73.054 61.629 ;
        RECT 72.726 55.121 72.772 61.911 ;
        RECT 65.964 61.883 72.726 61.957 ;
        RECT 66.332 61.515 73.1 61.583 ;
        RECT 72.68 55.167 72.726 61.957 ;
        RECT 65.918 61.929 72.68 62.003 ;
        RECT 66.378 61.469 73.146 61.537 ;
        RECT 72.634 55.213 72.68 62.003 ;
        RECT 65.872 61.975 72.634 62.049 ;
        RECT 66.424 61.423 73.192 61.491 ;
        RECT 72.588 55.259 72.634 62.049 ;
        RECT 65.826 62.021 72.588 62.095 ;
        RECT 66.47 61.377 73.238 61.445 ;
        RECT 72.542 55.305 72.588 62.095 ;
        RECT 65.78 62.067 72.542 62.141 ;
        RECT 66.516 61.331 73.284 61.399 ;
        RECT 72.496 55.351 72.542 62.141 ;
        RECT 65.734 62.113 72.496 62.187 ;
        RECT 66.562 61.285 73.33 61.353 ;
        RECT 72.45 55.397 72.496 62.187 ;
        RECT 65.688 62.159 72.45 62.233 ;
        RECT 66.608 61.239 73.376 61.307 ;
        RECT 72.404 55.443 72.45 62.233 ;
        RECT 65.642 62.205 72.404 62.279 ;
        RECT 66.654 61.193 73.422 61.261 ;
        RECT 72.358 55.489 72.404 62.279 ;
        RECT 65.596 62.251 72.358 62.325 ;
        RECT 66.7 61.147 73.468 61.215 ;
        RECT 72.312 55.535 72.358 62.325 ;
        RECT 65.55 62.297 72.312 62.371 ;
        RECT 66.746 61.101 73.514 61.169 ;
        RECT 72.266 55.581 72.312 62.371 ;
        RECT 65.504 62.343 72.266 62.417 ;
        RECT 66.792 61.055 73.56 61.123 ;
        RECT 72.22 55.627 72.266 62.417 ;
        RECT 65.458 62.389 72.22 62.463 ;
        RECT 66.838 61.009 73.606 61.077 ;
        RECT 72.174 55.673 72.22 62.463 ;
        RECT 65.412 62.435 72.174 62.509 ;
        RECT 66.884 60.963 73.652 61.031 ;
        RECT 72.128 55.719 72.174 62.509 ;
        RECT 65.366 62.481 72.128 62.555 ;
        RECT 66.93 60.917 73.698 60.985 ;
        RECT 72.082 55.765 72.128 62.555 ;
        RECT 65.32 62.527 72.082 62.601 ;
        RECT 66.976 60.871 73.744 60.939 ;
        RECT 72.036 55.811 72.082 62.601 ;
        RECT 65.274 62.573 72.036 62.647 ;
        RECT 67.022 60.825 73.79 60.893 ;
        RECT 71.99 55.857 72.036 62.647 ;
        RECT 65.228 62.619 71.99 62.693 ;
        RECT 67.068 60.779 73.836 60.847 ;
        RECT 71.944 55.903 71.99 62.693 ;
        RECT 65.182 62.665 71.944 62.739 ;
        RECT 67.114 60.733 73.882 60.801 ;
        RECT 71.898 55.949 71.944 62.739 ;
        RECT 65.136 62.711 71.898 62.785 ;
        RECT 67.16 60.687 73.928 60.755 ;
        RECT 71.852 55.995 71.898 62.785 ;
        RECT 65.09 62.757 71.852 62.831 ;
        RECT 67.206 60.641 73.974 60.709 ;
        RECT 71.806 56.041 71.852 62.831 ;
        RECT 65.044 62.803 71.806 62.877 ;
        RECT 67.252 60.595 74.02 60.663 ;
        RECT 71.76 56.087 71.806 62.877 ;
        RECT 64.998 62.849 71.76 62.923 ;
        RECT 67.298 60.549 74.066 60.617 ;
        RECT 71.714 56.133 71.76 62.923 ;
        RECT 64.952 62.895 71.714 62.969 ;
        RECT 67.344 60.503 74.112 60.571 ;
        RECT 71.668 56.179 71.714 62.969 ;
        RECT 64.906 62.941 71.668 63.015 ;
        RECT 67.39 60.457 74.158 60.525 ;
        RECT 71.622 56.225 71.668 63.015 ;
        RECT 64.86 62.987 71.622 63.061 ;
        RECT 67.436 60.411 74.204 60.479 ;
        RECT 71.576 56.271 71.622 63.061 ;
        RECT 64.814 63.033 71.576 63.107 ;
        RECT 67.482 60.365 74.25 60.433 ;
        RECT 71.53 56.317 71.576 63.107 ;
        RECT 64.768 63.079 71.53 63.153 ;
        RECT 67.528 60.319 74.296 60.387 ;
        RECT 71.484 56.363 71.53 63.153 ;
        RECT 64.722 63.125 71.484 63.199 ;
        RECT 67.574 60.273 74.342 60.341 ;
        RECT 71.438 56.409 71.484 63.199 ;
        RECT 64.676 63.171 71.438 63.245 ;
        RECT 67.62 60.227 74.388 60.295 ;
        RECT 71.392 56.455 71.438 63.245 ;
        RECT 64.63 63.217 71.392 63.291 ;
        RECT 67.666 60.181 74.434 60.249 ;
        RECT 71.346 56.501 71.392 63.291 ;
        RECT 64.584 63.263 71.346 63.337 ;
        RECT 67.712 60.135 74.48 60.203 ;
        RECT 71.3 56.547 71.346 63.337 ;
        RECT 64.538 63.309 71.3 63.383 ;
        RECT 67.758 60.089 74.526 60.157 ;
        RECT 71.254 56.593 71.3 63.383 ;
        RECT 64.492 63.355 71.254 63.429 ;
        RECT 67.804 60.043 74.572 60.111 ;
        RECT 71.208 56.639 71.254 63.429 ;
        RECT 64.446 63.401 71.208 63.475 ;
        RECT 67.85 59.997 74.618 60.065 ;
        RECT 71.162 56.685 71.208 63.475 ;
        RECT 64.4 63.447 71.162 63.521 ;
        RECT 67.896 59.951 74.664 60.019 ;
        RECT 71.116 56.731 71.162 63.521 ;
        RECT 64.354 63.493 71.116 63.567 ;
        RECT 67.942 59.905 74.71 59.973 ;
        RECT 71.07 56.777 71.116 63.567 ;
        RECT 64.308 63.539 71.07 63.613 ;
        RECT 67.988 59.859 74.756 59.927 ;
        RECT 71.024 56.823 71.07 63.613 ;
        RECT 64.262 63.585 71.024 63.659 ;
        RECT 68.034 59.813 74.802 59.881 ;
        RECT 70.978 56.869 71.024 63.659 ;
        RECT 64.216 63.631 70.978 63.705 ;
        RECT 68.08 59.767 74.848 59.835 ;
        RECT 70.932 56.915 70.978 63.705 ;
        RECT 64.17 63.677 70.932 63.751 ;
        RECT 68.126 59.721 80 59.8 ;
        RECT 70.886 56.961 70.932 63.751 ;
        RECT 64.124 63.723 70.886 63.797 ;
        RECT 68.172 59.675 80 59.8 ;
        RECT 70.84 57.007 70.886 63.797 ;
        RECT 64.078 63.769 70.84 63.843 ;
        RECT 68.218 59.629 80 59.8 ;
        RECT 70.794 57.053 70.84 63.843 ;
        RECT 64.032 63.815 70.794 63.889 ;
        RECT 68.264 59.583 80 59.8 ;
        RECT 70.748 57.099 70.794 63.889 ;
        RECT 63.986 63.861 70.748 63.935 ;
        RECT 68.31 59.537 80 59.8 ;
        RECT 70.702 57.145 70.748 63.935 ;
        RECT 63.94 63.907 70.702 63.981 ;
        RECT 68.356 59.491 80 59.8 ;
        RECT 70.656 57.191 70.702 63.981 ;
        RECT 63.894 63.953 70.656 64.027 ;
        RECT 68.402 59.445 80 59.8 ;
        RECT 70.61 57.237 70.656 64.027 ;
        RECT 63.848 63.999 70.61 64.073 ;
        RECT 68.448 59.399 80 59.8 ;
        RECT 70.564 57.283 70.61 64.073 ;
        RECT 63.802 64.045 70.564 64.119 ;
        RECT 68.494 59.353 80 59.8 ;
        RECT 70.518 57.329 70.564 64.119 ;
        RECT 63.756 64.091 70.518 64.165 ;
        RECT 68.54 59.307 80 59.8 ;
        RECT 70.472 57.375 70.518 64.165 ;
        RECT 63.71 64.137 70.472 64.211 ;
        RECT 68.586 59.261 80 59.8 ;
        RECT 70.426 57.421 70.472 64.211 ;
        RECT 63.664 64.183 70.426 64.257 ;
        RECT 68.632 59.215 80 59.8 ;
        RECT 70.38 57.467 70.426 64.257 ;
        RECT 63.618 64.229 70.38 64.303 ;
        RECT 68.678 59.169 80 59.8 ;
        RECT 70.334 57.513 70.38 64.303 ;
        RECT 63.572 64.275 70.334 64.349 ;
        RECT 68.724 59.123 80 59.8 ;
        RECT 70.288 57.559 70.334 64.349 ;
        RECT 63.526 64.321 70.288 64.395 ;
        RECT 68.77 59.077 80 59.8 ;
        RECT 70.242 57.605 70.288 64.395 ;
        RECT 63.48 64.367 70.242 64.441 ;
        RECT 68.816 59.031 80 59.8 ;
        RECT 70.196 57.651 70.242 64.441 ;
        RECT 63.434 64.413 70.196 64.487 ;
        RECT 68.862 58.985 80 59.8 ;
        RECT 70.15 57.697 70.196 64.487 ;
        RECT 63.388 64.459 70.15 64.533 ;
        RECT 68.908 58.939 80 59.8 ;
        RECT 70.104 57.743 70.15 64.533 ;
        RECT 63.342 64.505 70.104 64.579 ;
        RECT 68.954 58.893 80 59.8 ;
        RECT 70.058 57.789 70.104 64.579 ;
        RECT 63.296 64.551 70.058 64.625 ;
        RECT 69 58.847 80 59.8 ;
        RECT 70.012 57.835 70.058 64.625 ;
        RECT 63.25 64.597 70.012 64.671 ;
        RECT 69.046 58.801 80 59.8 ;
        RECT 69.966 57.881 70.012 64.671 ;
        RECT 63.204 64.643 69.966 64.717 ;
        RECT 69.092 58.755 80 59.8 ;
        RECT 69.92 57.927 69.966 64.717 ;
        RECT 63.158 64.689 69.92 64.763 ;
        RECT 69.138 58.709 80 59.8 ;
        RECT 69.874 57.973 69.92 64.763 ;
        RECT 63.112 64.735 69.874 64.809 ;
        RECT 69.184 58.663 80 59.8 ;
        RECT 69.828 58.019 69.874 64.809 ;
        RECT 63.066 64.781 69.828 64.855 ;
        RECT 69.23 58.617 80 59.8 ;
        RECT 69.782 58.065 69.828 64.855 ;
        RECT 63.02 64.827 69.782 64.901 ;
        RECT 69.276 58.571 80 59.8 ;
        RECT 69.736 58.111 69.782 64.901 ;
        RECT 62.974 64.873 69.736 64.947 ;
        RECT 69.322 58.525 80 59.8 ;
        RECT 69.69 58.157 69.736 64.947 ;
        RECT 62.928 64.919 69.69 64.993 ;
        RECT 69.368 58.479 80 59.8 ;
        RECT 69.644 58.203 69.69 64.993 ;
        RECT 62.882 64.965 69.644 65.039 ;
        RECT 69.414 58.433 80 59.8 ;
        RECT 69.598 58.249 69.644 65.039 ;
        RECT 62.836 65.011 69.598 65.085 ;
        RECT 69.46 58.387 80 59.8 ;
        RECT 69.552 58.295 69.598 65.085 ;
        RECT 62.79 65.057 69.552 65.131 ;
        RECT 69.506 58.341 80 59.8 ;
        RECT 62.744 65.103 69.506 65.177 ;
        RECT 62.698 65.149 69.46 65.223 ;
        RECT 62.652 65.195 69.414 65.269 ;
        RECT 62.606 65.241 69.368 65.315 ;
        RECT 62.56 65.287 69.322 65.361 ;
        RECT 62.514 65.333 69.276 65.407 ;
        RECT 62.468 65.379 69.23 65.453 ;
        RECT 62.422 65.425 69.184 65.499 ;
        RECT 62.376 65.471 69.138 65.545 ;
        RECT 62.33 65.517 69.092 65.591 ;
        RECT 62.284 65.563 69.046 65.637 ;
        RECT 62.238 65.609 69 65.683 ;
        RECT 62.192 65.655 68.954 65.729 ;
        RECT 62.146 65.701 68.908 65.775 ;
        RECT 62.1 65.747 68.862 65.821 ;
        RECT 62.054 65.793 68.816 65.867 ;
        RECT 62.008 65.839 68.77 65.913 ;
        RECT 61.962 65.885 68.724 65.959 ;
        RECT 61.916 65.931 68.678 66.005 ;
        RECT 61.87 65.977 68.632 66.051 ;
        RECT 61.824 66.023 68.586 66.097 ;
        RECT 61.778 66.069 68.54 66.143 ;
        RECT 61.732 66.115 68.494 66.189 ;
        RECT 61.686 66.161 68.448 66.235 ;
        RECT 61.64 66.207 68.402 66.281 ;
        RECT 61.594 66.253 68.356 66.327 ;
        RECT 61.548 66.299 68.31 66.373 ;
        RECT 61.502 66.345 68.264 66.419 ;
        RECT 61.456 66.391 68.218 66.465 ;
        RECT 61.41 66.437 68.172 66.511 ;
        RECT 61.364 66.483 68.126 66.557 ;
        RECT 61.318 66.529 68.08 66.603 ;
        RECT 61.272 66.575 68.034 66.649 ;
        RECT 61.226 66.621 67.988 66.695 ;
        RECT 61.18 66.667 67.942 66.741 ;
        RECT 61.134 66.713 67.896 66.787 ;
        RECT 61.088 66.759 67.85 66.833 ;
        RECT 61.042 66.805 67.804 66.879 ;
        RECT 60.996 66.851 67.758 66.925 ;
        RECT 60.95 66.897 67.712 66.971 ;
        RECT 60.904 66.943 67.666 67.017 ;
        RECT 60.858 66.989 67.62 67.063 ;
        RECT 60.812 67.035 67.574 67.109 ;
        RECT 60.766 67.081 67.528 67.155 ;
        RECT 60.72 67.127 67.482 67.201 ;
        RECT 60.674 67.173 67.436 67.247 ;
        RECT 60.628 67.219 67.39 67.293 ;
        RECT 60.582 67.265 67.344 67.339 ;
        RECT 60.536 67.311 67.298 67.385 ;
        RECT 60.49 67.357 67.252 67.431 ;
        RECT 60.444 67.403 67.206 67.477 ;
        RECT 60.398 67.449 67.16 67.523 ;
        RECT 60.352 67.495 67.114 67.569 ;
        RECT 60.306 67.541 67.068 67.615 ;
        RECT 60.26 67.587 67.022 67.661 ;
        RECT 60.214 67.633 66.976 67.707 ;
        RECT 60.168 67.679 66.93 67.753 ;
        RECT 60.122 67.725 66.884 67.799 ;
        RECT 60.076 67.771 66.838 67.845 ;
        RECT 60.03 67.817 66.792 67.891 ;
        RECT 59.984 67.863 66.746 67.937 ;
        RECT 59.938 67.909 66.7 67.983 ;
        RECT 59.892 67.955 66.654 68.029 ;
        RECT 59.846 68.001 66.608 68.075 ;
        RECT 59.784 68.078 66.562 68.121 ;
        RECT 59.8 68.047 66.562 68.121 ;
        RECT 59.738 68.109 66.516 68.167 ;
        RECT 59.692 68.155 66.47 68.213 ;
        RECT 59.646 68.201 66.424 68.259 ;
        RECT 59.6 68.247 66.378 68.305 ;
        RECT 59.554 68.293 66.332 68.351 ;
        RECT 59.508 68.339 66.286 68.397 ;
        RECT 59.462 68.385 66.24 68.443 ;
        RECT 59.416 68.431 66.194 68.489 ;
        RECT 59.37 68.477 66.148 68.535 ;
        RECT 59.324 68.523 66.102 68.581 ;
        RECT 59.278 68.569 66.056 68.627 ;
        RECT 59.232 68.615 66.01 68.673 ;
        RECT 59.186 68.661 65.964 68.719 ;
        RECT 59.14 68.707 65.918 68.765 ;
        RECT 59.094 68.753 65.872 68.811 ;
        RECT 59.048 68.799 65.826 68.857 ;
        RECT 59.002 68.845 65.78 68.903 ;
        RECT 58.956 68.891 65.734 68.949 ;
        RECT 58.91 68.937 65.688 68.995 ;
        RECT 58.864 68.983 65.642 69.041 ;
        RECT 58.818 69.029 65.596 69.087 ;
        RECT 58.772 69.075 65.55 69.133 ;
        RECT 58.726 69.121 65.504 69.179 ;
        RECT 58.68 69.167 65.458 69.225 ;
        RECT 58.634 69.213 65.412 69.271 ;
        RECT 58.588 69.259 65.366 69.317 ;
        RECT 58.542 69.305 65.32 69.363 ;
        RECT 58.496 69.351 65.274 69.409 ;
        RECT 58.45 69.397 65.228 69.455 ;
        RECT 58.404 69.443 65.182 69.501 ;
        RECT 58.358 69.489 65.136 69.547 ;
        RECT 58.312 69.535 65.09 69.593 ;
        RECT 58.266 69.581 65.044 69.639 ;
        RECT 58.22 69.627 64.998 69.685 ;
        RECT 58.174 69.673 64.952 69.731 ;
        RECT 58.128 69.719 64.906 69.777 ;
        RECT 58.082 69.765 64.86 69.823 ;
        RECT 58.036 69.811 64.814 69.869 ;
        RECT 57.99 69.857 64.768 69.915 ;
        RECT 57.944 69.903 64.722 69.961 ;
        RECT 57.898 69.949 64.676 70.007 ;
        RECT 57.852 69.995 64.63 70.053 ;
        RECT 57.806 70.041 64.584 70.099 ;
        RECT 57.76 70.087 64.538 70.145 ;
        RECT 57.714 70.133 64.492 70.191 ;
        RECT 57.668 70.179 64.446 70.237 ;
        RECT 57.622 70.225 64.4 70.283 ;
        RECT 57.576 70.271 64.354 70.329 ;
        RECT 57.53 70.317 64.308 70.375 ;
        RECT 57.484 70.363 64.262 70.421 ;
        RECT 57.438 70.409 64.216 70.467 ;
        RECT 57.392 70.455 64.17 70.513 ;
        RECT 57.346 70.501 64.124 70.559 ;
        RECT 57.3 70.547 64.078 70.605 ;
        RECT 57.254 70.593 64.032 70.651 ;
        RECT 57.208 70.639 63.986 70.697 ;
        RECT 57.162 70.685 63.94 70.743 ;
        RECT 57.116 70.731 63.894 70.789 ;
        RECT 57.07 70.777 63.848 70.835 ;
        RECT 57.024 70.823 63.802 70.881 ;
        RECT 56.978 70.869 63.756 70.927 ;
        RECT 56.932 70.915 63.71 70.973 ;
        RECT 56.886 70.961 63.664 71.019 ;
        RECT 56.84 71.007 63.618 71.065 ;
        RECT 56.794 71.053 63.572 71.111 ;
        RECT 56.748 71.099 63.526 71.157 ;
        RECT 56.702 71.145 63.48 71.203 ;
        RECT 56.656 71.191 63.434 71.249 ;
        RECT 56.61 71.237 63.388 71.295 ;
        RECT 56.564 71.283 63.342 71.341 ;
        RECT 56.518 71.329 63.296 71.387 ;
        RECT 56.472 71.375 63.25 71.433 ;
        RECT 56.426 71.421 63.204 71.479 ;
        RECT 56.38 71.467 63.158 71.525 ;
        RECT 56.334 71.513 63.112 71.571 ;
        RECT 56.288 71.559 63.066 71.617 ;
        RECT 56.242 71.605 63.02 71.663 ;
        RECT 56.196 71.651 62.974 71.709 ;
        RECT 56.15 71.697 62.928 71.755 ;
        RECT 56.104 71.743 62.882 71.801 ;
        RECT 56.058 71.789 62.836 71.847 ;
        RECT 56.012 71.835 62.79 71.893 ;
        RECT 55.966 71.881 62.744 71.939 ;
        RECT 55.92 71.927 62.698 71.985 ;
        RECT 55.874 71.973 62.652 72.031 ;
        RECT 55.828 72.019 62.606 72.077 ;
        RECT 55.782 72.065 62.56 72.123 ;
        RECT 55.736 72.111 62.514 72.169 ;
        RECT 55.69 72.157 62.468 72.215 ;
        RECT 55.644 72.203 62.422 72.261 ;
        RECT 55.598 72.249 62.376 72.307 ;
        RECT 55.552 72.295 62.33 72.353 ;
        RECT 55.506 72.341 62.284 72.399 ;
        RECT 55.46 72.387 62.238 72.445 ;
        RECT 55.414 72.433 62.192 72.491 ;
        RECT 55.368 72.479 62.146 72.537 ;
        RECT 55.322 72.525 62.1 72.583 ;
        RECT 55.276 72.571 62.054 72.629 ;
        RECT 55.23 72.617 62.008 72.675 ;
        RECT 55.184 72.663 61.962 72.721 ;
        RECT 55.138 72.709 61.916 72.767 ;
        RECT 55.092 72.755 61.87 72.813 ;
        RECT 55.046 72.801 61.824 72.859 ;
        RECT 55 72.847 61.778 72.905 ;
        RECT 55 72.847 61.732 72.951 ;
        RECT 55 72.847 61.686 72.997 ;
        RECT 55 72.847 61.64 73.043 ;
        RECT 55 72.847 61.594 73.089 ;
        RECT 55 72.847 61.548 73.135 ;
        RECT 55 72.847 61.502 73.181 ;
        RECT 55 72.847 61.456 73.227 ;
        RECT 55 72.847 61.41 73.273 ;
        RECT 55 72.847 61.364 73.319 ;
        RECT 55 72.847 61.318 73.365 ;
        RECT 55 72.847 61.272 73.411 ;
        RECT 55 72.847 61.226 73.457 ;
        RECT 55 72.847 61.18 73.503 ;
        RECT 55 72.847 61.134 73.549 ;
        RECT 55 72.847 61.088 73.595 ;
        RECT 55 72.847 61.042 73.641 ;
        RECT 55 72.847 60.996 73.687 ;
        RECT 55 72.847 60.95 73.733 ;
        RECT 55 72.847 60.904 73.779 ;
        RECT 55 72.847 60.858 73.825 ;
        RECT 55 72.847 60.812 73.871 ;
        RECT 55 72.847 60.766 73.917 ;
        RECT 55 72.847 60.72 73.963 ;
        RECT 55 72.847 60.674 74.009 ;
        RECT 55 72.847 60.628 74.055 ;
        RECT 55 72.847 60.582 74.101 ;
        RECT 55 72.847 60.536 74.147 ;
        RECT 55 72.847 60.49 74.193 ;
        RECT 55 72.847 60.444 74.239 ;
        RECT 55 72.847 60.398 74.285 ;
        RECT 55 72.847 60.352 74.331 ;
        RECT 55 72.847 60.306 74.377 ;
        RECT 55 72.847 60.26 74.423 ;
        RECT 55 72.847 60.214 74.469 ;
        RECT 55 72.847 60.168 74.515 ;
        RECT 55 72.847 60.122 74.561 ;
        RECT 55 72.847 60.076 74.607 ;
        RECT 55 72.847 60.03 74.653 ;
        RECT 55 72.847 59.984 74.699 ;
        RECT 55 72.847 59.938 74.745 ;
        RECT 55 72.847 59.892 74.791 ;
        RECT 55 72.847 59.846 74.837 ;
        RECT 55 72.847 59.8 80 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 62.59 30.2 80 35 ;
        RECT 57.77 34.997 64.58 35.006 ;
        RECT 57.77 34.997 64.568 35.035 ;
        RECT 55.838 36.929 62.59 37.008 ;
        RECT 55.884 36.883 62.636 36.967 ;
        RECT 62.554 30.218 62.59 37.008 ;
        RECT 55.792 36.975 62.554 37.049 ;
        RECT 55.93 36.837 62.682 36.921 ;
        RECT 62.508 30.259 62.554 37.049 ;
        RECT 55.746 37.021 62.508 37.095 ;
        RECT 55.976 36.791 62.728 36.875 ;
        RECT 62.462 30.305 62.508 37.095 ;
        RECT 55.7 37.067 62.462 37.141 ;
        RECT 56.022 36.745 62.774 36.829 ;
        RECT 62.416 30.351 62.462 37.141 ;
        RECT 55.654 37.113 62.416 37.187 ;
        RECT 56.068 36.699 62.82 36.783 ;
        RECT 62.37 30.397 62.416 37.187 ;
        RECT 55.608 37.159 62.37 37.233 ;
        RECT 56.114 36.653 62.866 36.737 ;
        RECT 62.324 30.443 62.37 37.233 ;
        RECT 55.562 37.205 62.324 37.279 ;
        RECT 56.16 36.607 62.912 36.691 ;
        RECT 62.278 30.489 62.324 37.279 ;
        RECT 55.516 37.251 62.278 37.325 ;
        RECT 56.206 36.561 62.958 36.645 ;
        RECT 62.232 30.535 62.278 37.325 ;
        RECT 55.47 37.297 62.232 37.371 ;
        RECT 56.252 36.515 63.004 36.599 ;
        RECT 62.186 30.581 62.232 37.371 ;
        RECT 55.424 37.343 62.186 37.417 ;
        RECT 56.298 36.469 63.05 36.553 ;
        RECT 62.14 30.627 62.186 37.417 ;
        RECT 55.378 37.389 62.14 37.463 ;
        RECT 56.344 36.423 63.096 36.507 ;
        RECT 62.094 30.673 62.14 37.463 ;
        RECT 55.332 37.435 62.094 37.509 ;
        RECT 56.39 36.377 63.142 36.461 ;
        RECT 62.048 30.719 62.094 37.509 ;
        RECT 55.286 37.481 62.048 37.555 ;
        RECT 56.436 36.331 63.188 36.415 ;
        RECT 62.002 30.765 62.048 37.555 ;
        RECT 55.24 37.527 62.002 37.601 ;
        RECT 56.482 36.285 63.234 36.369 ;
        RECT 61.956 30.811 62.002 37.601 ;
        RECT 55.194 37.573 61.956 37.647 ;
        RECT 56.528 36.239 63.28 36.323 ;
        RECT 61.91 30.857 61.956 37.647 ;
        RECT 55.148 37.619 61.91 37.693 ;
        RECT 56.574 36.193 63.326 36.277 ;
        RECT 61.864 30.903 61.91 37.693 ;
        RECT 55.102 37.665 61.864 37.739 ;
        RECT 56.62 36.147 63.372 36.231 ;
        RECT 61.818 30.949 61.864 37.739 ;
        RECT 55.056 37.711 61.818 37.785 ;
        RECT 56.666 36.101 63.418 36.185 ;
        RECT 61.772 30.995 61.818 37.785 ;
        RECT 55.01 37.757 61.772 37.831 ;
        RECT 56.712 36.055 63.464 36.139 ;
        RECT 61.726 31.041 61.772 37.831 ;
        RECT 54.964 37.803 61.726 37.877 ;
        RECT 56.758 36.009 63.51 36.093 ;
        RECT 61.68 31.087 61.726 37.877 ;
        RECT 54.918 37.849 61.68 37.923 ;
        RECT 56.804 35.963 63.556 36.047 ;
        RECT 61.634 31.133 61.68 37.923 ;
        RECT 54.872 37.895 61.634 37.969 ;
        RECT 56.85 35.917 63.602 36.001 ;
        RECT 61.588 31.179 61.634 37.969 ;
        RECT 54.826 37.941 61.588 38.015 ;
        RECT 56.896 35.871 63.648 35.955 ;
        RECT 61.542 31.225 61.588 38.015 ;
        RECT 54.78 37.987 61.542 38.061 ;
        RECT 56.942 35.825 63.694 35.909 ;
        RECT 61.496 31.271 61.542 38.061 ;
        RECT 54.734 38.033 61.496 38.107 ;
        RECT 56.988 35.779 63.74 35.863 ;
        RECT 61.45 31.317 61.496 38.107 ;
        RECT 54.688 38.079 61.45 38.153 ;
        RECT 57.034 35.733 63.786 35.817 ;
        RECT 61.404 31.363 61.45 38.153 ;
        RECT 54.642 38.125 61.404 38.199 ;
        RECT 57.08 35.687 63.832 35.771 ;
        RECT 61.358 31.409 61.404 38.199 ;
        RECT 54.596 38.171 61.358 38.245 ;
        RECT 57.126 35.641 63.878 35.725 ;
        RECT 61.312 31.455 61.358 38.245 ;
        RECT 54.55 38.217 61.312 38.291 ;
        RECT 57.172 35.595 63.924 35.679 ;
        RECT 61.266 31.501 61.312 38.291 ;
        RECT 54.504 38.263 61.266 38.337 ;
        RECT 57.218 35.549 63.97 35.633 ;
        RECT 61.22 31.547 61.266 38.337 ;
        RECT 54.458 38.309 61.22 38.383 ;
        RECT 57.264 35.503 64.016 35.587 ;
        RECT 61.174 31.593 61.22 38.383 ;
        RECT 54.412 38.355 61.174 38.429 ;
        RECT 57.31 35.457 64.062 35.541 ;
        RECT 61.128 31.639 61.174 38.429 ;
        RECT 54.366 38.401 61.128 38.475 ;
        RECT 57.356 35.411 64.108 35.495 ;
        RECT 61.082 31.685 61.128 38.475 ;
        RECT 54.32 38.447 61.082 38.521 ;
        RECT 57.402 35.365 64.154 35.449 ;
        RECT 61.036 31.731 61.082 38.521 ;
        RECT 54.274 38.493 61.036 38.567 ;
        RECT 57.448 35.319 64.2 35.403 ;
        RECT 60.99 31.777 61.036 38.567 ;
        RECT 54.228 38.539 60.99 38.613 ;
        RECT 57.494 35.273 64.246 35.357 ;
        RECT 60.944 31.823 60.99 38.613 ;
        RECT 54.182 38.585 60.944 38.659 ;
        RECT 57.54 35.227 64.292 35.311 ;
        RECT 60.898 31.869 60.944 38.659 ;
        RECT 54.136 38.631 60.898 38.705 ;
        RECT 57.586 35.181 64.338 35.265 ;
        RECT 60.852 31.915 60.898 38.705 ;
        RECT 54.09 38.677 60.852 38.751 ;
        RECT 57.632 35.135 64.384 35.219 ;
        RECT 60.806 31.961 60.852 38.751 ;
        RECT 54.044 38.723 60.806 38.797 ;
        RECT 57.678 35.089 64.43 35.173 ;
        RECT 60.76 32.007 60.806 38.797 ;
        RECT 53.998 38.769 60.76 38.843 ;
        RECT 57.724 35.043 64.476 35.127 ;
        RECT 60.714 32.053 60.76 38.843 ;
        RECT 53.952 38.815 60.714 38.889 ;
        RECT 57.77 34.997 64.522 35.081 ;
        RECT 60.668 32.099 60.714 38.889 ;
        RECT 53.906 38.861 60.668 38.935 ;
        RECT 57.816 34.951 80 35 ;
        RECT 60.622 32.145 60.668 38.935 ;
        RECT 53.86 38.907 60.622 38.981 ;
        RECT 57.862 34.905 80 35 ;
        RECT 60.576 32.191 60.622 38.981 ;
        RECT 53.814 38.953 60.576 39.027 ;
        RECT 57.908 34.859 80 35 ;
        RECT 60.53 32.237 60.576 39.027 ;
        RECT 53.768 38.999 60.53 39.073 ;
        RECT 57.954 34.813 80 35 ;
        RECT 60.484 32.283 60.53 39.073 ;
        RECT 53.722 39.045 60.484 39.119 ;
        RECT 58 34.767 80 35 ;
        RECT 60.438 32.329 60.484 39.119 ;
        RECT 53.676 39.091 60.438 39.165 ;
        RECT 58.046 34.721 80 35 ;
        RECT 60.392 32.375 60.438 39.165 ;
        RECT 53.63 39.137 60.392 39.211 ;
        RECT 58.092 34.675 80 35 ;
        RECT 60.346 32.421 60.392 39.211 ;
        RECT 53.584 39.183 60.346 39.257 ;
        RECT 58.138 34.629 80 35 ;
        RECT 60.3 32.467 60.346 39.257 ;
        RECT 53.538 39.229 60.3 39.303 ;
        RECT 58.184 34.583 80 35 ;
        RECT 60.254 32.513 60.3 39.303 ;
        RECT 53.492 39.275 60.254 39.349 ;
        RECT 58.23 34.537 80 35 ;
        RECT 60.208 32.559 60.254 39.349 ;
        RECT 53.446 39.321 60.208 39.395 ;
        RECT 58.276 34.491 80 35 ;
        RECT 60.162 32.605 60.208 39.395 ;
        RECT 53.4 39.367 60.162 39.441 ;
        RECT 58.322 34.445 80 35 ;
        RECT 60.116 32.651 60.162 39.441 ;
        RECT 53.354 39.413 60.116 39.487 ;
        RECT 58.368 34.399 80 35 ;
        RECT 60.07 32.697 60.116 39.487 ;
        RECT 53.308 39.459 60.07 39.533 ;
        RECT 58.414 34.353 80 35 ;
        RECT 60.024 32.743 60.07 39.533 ;
        RECT 53.262 39.505 60.024 39.579 ;
        RECT 58.46 34.307 80 35 ;
        RECT 59.978 32.789 60.024 39.579 ;
        RECT 53.216 39.551 59.978 39.625 ;
        RECT 58.506 34.261 80 35 ;
        RECT 59.932 32.835 59.978 39.625 ;
        RECT 53.17 39.597 59.932 39.671 ;
        RECT 58.552 34.215 80 35 ;
        RECT 59.886 32.881 59.932 39.671 ;
        RECT 53.124 39.643 59.886 39.717 ;
        RECT 58.598 34.169 80 35 ;
        RECT 59.84 32.927 59.886 39.717 ;
        RECT 53.078 39.689 59.84 39.763 ;
        RECT 58.644 34.123 80 35 ;
        RECT 59.794 32.973 59.84 39.763 ;
        RECT 53.032 39.735 59.794 39.809 ;
        RECT 58.69 34.077 80 35 ;
        RECT 59.748 33.019 59.794 39.809 ;
        RECT 52.986 39.781 59.748 39.855 ;
        RECT 58.736 34.031 80 35 ;
        RECT 59.702 33.065 59.748 39.855 ;
        RECT 52.94 39.827 59.702 39.901 ;
        RECT 58.782 33.985 80 35 ;
        RECT 59.656 33.111 59.702 39.901 ;
        RECT 52.894 39.873 59.656 39.947 ;
        RECT 58.828 33.939 80 35 ;
        RECT 59.61 33.157 59.656 39.947 ;
        RECT 52.848 39.919 59.61 39.993 ;
        RECT 58.874 33.893 80 35 ;
        RECT 59.564 33.203 59.61 39.993 ;
        RECT 52.802 39.965 59.564 40.039 ;
        RECT 58.92 33.847 80 35 ;
        RECT 59.518 33.249 59.564 40.039 ;
        RECT 52.756 40.011 59.518 40.085 ;
        RECT 58.966 33.801 80 35 ;
        RECT 59.472 33.295 59.518 40.085 ;
        RECT 52.71 40.057 59.472 40.131 ;
        RECT 59.012 33.755 80 35 ;
        RECT 59.426 33.341 59.472 40.131 ;
        RECT 52.664 40.103 59.426 40.177 ;
        RECT 59.058 33.709 80 35 ;
        RECT 59.38 33.387 59.426 40.177 ;
        RECT 52.618 40.149 59.38 40.223 ;
        RECT 59.104 33.663 80 35 ;
        RECT 59.334 33.433 59.38 40.223 ;
        RECT 52.572 40.195 59.334 40.269 ;
        RECT 59.15 33.617 80 35 ;
        RECT 59.288 33.479 59.334 40.269 ;
        RECT 52.526 40.241 59.288 40.315 ;
        RECT 59.196 33.571 80 35 ;
        RECT 59.242 33.525 59.288 40.315 ;
        RECT 52.48 40.287 59.242 40.361 ;
        RECT 52.434 40.333 59.196 40.407 ;
        RECT 52.388 40.379 59.15 40.453 ;
        RECT 52.342 40.425 59.104 40.499 ;
        RECT 52.296 40.471 59.058 40.545 ;
        RECT 52.25 40.517 59.012 40.591 ;
        RECT 52.204 40.563 58.966 40.637 ;
        RECT 52.158 40.609 58.92 40.683 ;
        RECT 52.112 40.655 58.874 40.729 ;
        RECT 52.066 40.701 58.828 40.775 ;
        RECT 52.02 40.747 58.782 40.821 ;
        RECT 51.974 40.793 58.736 40.867 ;
        RECT 51.928 40.839 58.69 40.913 ;
        RECT 51.882 40.885 58.644 40.959 ;
        RECT 51.836 40.931 58.598 41.005 ;
        RECT 51.79 40.977 58.552 41.051 ;
        RECT 51.744 41.023 58.506 41.097 ;
        RECT 51.698 41.069 58.46 41.143 ;
        RECT 51.652 41.115 58.414 41.189 ;
        RECT 51.606 41.161 58.368 41.235 ;
        RECT 51.56 41.207 58.322 41.281 ;
        RECT 51.514 41.253 58.276 41.327 ;
        RECT 51.468 41.299 58.23 41.373 ;
        RECT 51.422 41.345 58.184 41.419 ;
        RECT 51.376 41.391 58.138 41.465 ;
        RECT 51.33 41.437 58.092 41.511 ;
        RECT 51.284 41.483 58.046 41.557 ;
        RECT 51.238 41.529 58 41.603 ;
        RECT 51.192 41.575 57.954 41.649 ;
        RECT 51.146 41.621 57.908 41.695 ;
        RECT 51.1 41.667 57.862 41.741 ;
        RECT 51.054 41.713 57.816 41.787 ;
        RECT 51.008 41.759 57.77 41.833 ;
        RECT 50.962 41.805 57.724 41.879 ;
        RECT 50.916 41.851 57.678 41.925 ;
        RECT 50.87 41.897 57.632 41.971 ;
        RECT 50.824 41.943 57.586 42.017 ;
        RECT 50.778 41.989 57.54 42.063 ;
        RECT 50.732 42.035 57.494 42.109 ;
        RECT 50.686 42.081 57.448 42.155 ;
        RECT 50.64 42.127 57.402 42.201 ;
        RECT 50.594 42.173 57.356 42.247 ;
        RECT 50.548 42.219 57.31 42.293 ;
        RECT 50.502 42.265 57.264 42.339 ;
        RECT 50.456 42.311 57.218 42.385 ;
        RECT 50.41 42.357 57.172 42.431 ;
        RECT 50.364 42.403 57.126 42.477 ;
        RECT 50.318 42.449 57.08 42.523 ;
        RECT 50.272 42.495 57.034 42.569 ;
        RECT 50.226 42.541 56.988 42.615 ;
        RECT 50.18 42.587 56.942 42.661 ;
        RECT 50.134 42.633 56.896 42.707 ;
        RECT 50.088 42.679 56.85 42.753 ;
        RECT 50.042 42.725 56.804 42.799 ;
        RECT 49.996 42.771 56.758 42.845 ;
        RECT 49.95 42.817 56.712 42.891 ;
        RECT 49.904 42.863 56.666 42.937 ;
        RECT 49.858 42.909 56.62 42.983 ;
        RECT 49.812 42.955 56.574 43.029 ;
        RECT 49.766 43.001 56.528 43.075 ;
        RECT 49.72 43.047 56.482 43.121 ;
        RECT 49.674 43.093 56.436 43.167 ;
        RECT 49.628 43.139 56.39 43.213 ;
        RECT 49.582 43.185 56.344 43.259 ;
        RECT 49.536 43.231 56.298 43.305 ;
        RECT 49.49 43.277 56.252 43.351 ;
        RECT 49.444 43.323 56.206 43.397 ;
        RECT 49.398 43.369 56.16 43.443 ;
        RECT 49.352 43.415 56.114 43.489 ;
        RECT 49.306 43.461 56.068 43.535 ;
        RECT 49.26 43.507 56.022 43.581 ;
        RECT 49.214 43.553 55.976 43.627 ;
        RECT 49.168 43.599 55.93 43.673 ;
        RECT 49.122 43.645 55.884 43.719 ;
        RECT 49.076 43.691 55.838 43.765 ;
        RECT 49.03 43.737 55.792 43.811 ;
        RECT 48.984 43.783 55.746 43.857 ;
        RECT 48.938 43.829 55.7 43.903 ;
        RECT 48.892 43.875 55.654 43.949 ;
        RECT 48.846 43.921 55.608 43.995 ;
        RECT 48.8 43.967 55.562 44.041 ;
        RECT 48.754 44.013 55.516 44.087 ;
        RECT 48.708 44.059 55.47 44.133 ;
        RECT 48.662 44.105 55.424 44.179 ;
        RECT 48.616 44.151 55.378 44.225 ;
        RECT 48.57 44.197 55.332 44.271 ;
        RECT 48.524 44.243 55.286 44.317 ;
        RECT 48.478 44.289 55.24 44.363 ;
        RECT 48.432 44.335 55.194 44.409 ;
        RECT 48.386 44.381 55.148 44.455 ;
        RECT 48.34 44.427 55.102 44.501 ;
        RECT 48.294 44.473 55.056 44.547 ;
        RECT 48.248 44.519 55.01 44.593 ;
        RECT 48.202 44.565 54.964 44.639 ;
        RECT 48.156 44.611 54.918 44.685 ;
        RECT 48.11 44.657 54.872 44.731 ;
        RECT 48.064 44.703 54.826 44.777 ;
        RECT 48.018 44.749 54.78 44.823 ;
        RECT 47.972 44.795 54.734 44.869 ;
        RECT 47.926 44.841 54.688 44.915 ;
        RECT 47.88 44.887 54.642 44.961 ;
        RECT 47.834 44.933 54.596 45.007 ;
        RECT 47.788 44.979 54.55 45.053 ;
        RECT 47.742 45.025 54.504 45.099 ;
        RECT 47.696 45.071 54.458 45.145 ;
        RECT 47.65 45.117 54.412 45.191 ;
        RECT 47.604 45.163 54.366 45.237 ;
        RECT 47.558 45.209 54.32 45.283 ;
        RECT 47.512 45.255 54.274 45.329 ;
        RECT 47.466 45.301 54.228 45.375 ;
        RECT 47.42 45.347 54.182 45.421 ;
        RECT 47.374 45.393 54.136 45.467 ;
        RECT 47.328 45.439 54.09 45.513 ;
        RECT 47.282 45.485 54.044 45.559 ;
        RECT 47.236 45.531 53.998 45.605 ;
        RECT 47.19 45.577 53.952 45.651 ;
        RECT 47.144 45.623 53.906 45.697 ;
        RECT 47.098 45.669 53.86 45.743 ;
        RECT 47.052 45.715 53.814 45.789 ;
        RECT 47.006 45.761 53.768 45.835 ;
        RECT 46.96 45.807 53.722 45.881 ;
        RECT 46.914 45.853 53.676 45.927 ;
        RECT 46.868 45.899 53.63 45.973 ;
        RECT 46.822 45.945 53.584 46.019 ;
        RECT 46.776 45.991 53.538 46.065 ;
        RECT 46.73 46.037 53.492 46.111 ;
        RECT 46.684 46.083 53.446 46.157 ;
        RECT 46.638 46.129 53.4 46.203 ;
        RECT 46.592 46.175 53.354 46.249 ;
        RECT 46.546 46.221 53.308 46.295 ;
        RECT 46.5 46.267 53.262 46.341 ;
        RECT 46.454 46.313 53.216 46.387 ;
        RECT 46.408 46.359 53.17 46.433 ;
        RECT 46.362 46.405 53.124 46.479 ;
        RECT 46.316 46.451 53.078 46.525 ;
        RECT 46.27 46.497 53.032 46.571 ;
        RECT 46.224 46.543 52.986 46.617 ;
        RECT 46.178 46.589 52.94 46.663 ;
        RECT 46.132 46.635 52.894 46.709 ;
        RECT 46.086 46.681 52.848 46.755 ;
        RECT 46.04 46.727 52.802 46.801 ;
        RECT 45.994 46.773 52.756 46.847 ;
        RECT 45.948 46.819 52.71 46.893 ;
        RECT 45.902 46.865 52.664 46.939 ;
        RECT 45.856 46.911 52.618 46.985 ;
        RECT 45.81 46.957 52.572 47.031 ;
        RECT 45.764 47.003 52.526 47.077 ;
        RECT 45.718 47.049 52.48 47.123 ;
        RECT 45.672 47.095 52.434 47.169 ;
        RECT 45.626 47.141 52.388 47.215 ;
        RECT 45.58 47.187 52.342 47.261 ;
        RECT 45.534 47.233 52.296 47.307 ;
        RECT 45.488 47.279 52.25 47.353 ;
        RECT 45.442 47.325 52.204 47.399 ;
        RECT 45.396 47.371 52.158 47.445 ;
        RECT 45.35 47.417 52.112 47.491 ;
        RECT 45.304 47.463 52.066 47.537 ;
        RECT 45.258 47.509 52.02 47.583 ;
        RECT 45.212 47.555 51.974 47.629 ;
        RECT 45.166 47.601 51.928 47.675 ;
        RECT 45.12 47.647 51.882 47.721 ;
        RECT 45.074 47.693 51.836 47.767 ;
        RECT 45.028 47.739 51.79 47.813 ;
        RECT 44.982 47.785 51.744 47.859 ;
        RECT 44.936 47.831 51.698 47.905 ;
        RECT 44.89 47.877 51.652 47.951 ;
        RECT 44.844 47.923 51.606 47.997 ;
        RECT 44.798 47.969 51.56 48.043 ;
        RECT 44.752 48.015 51.514 48.089 ;
        RECT 44.706 48.061 51.468 48.135 ;
        RECT 44.66 48.107 51.422 48.181 ;
        RECT 44.614 48.153 51.376 48.227 ;
        RECT 44.568 48.199 51.33 48.273 ;
        RECT 44.522 48.245 51.284 48.319 ;
        RECT 44.476 48.291 51.238 48.365 ;
        RECT 44.43 48.337 51.192 48.411 ;
        RECT 44.384 48.383 51.146 48.457 ;
        RECT 44.338 48.429 51.1 48.503 ;
        RECT 44.292 48.475 51.054 48.549 ;
        RECT 44.246 48.521 51.008 48.595 ;
        RECT 44.2 48.567 50.962 48.641 ;
        RECT 44.154 48.613 50.916 48.687 ;
        RECT 44.108 48.659 50.87 48.733 ;
        RECT 44.062 48.705 50.824 48.779 ;
        RECT 44.016 48.751 50.778 48.825 ;
        RECT 43.97 48.797 50.732 48.871 ;
        RECT 43.924 48.843 50.686 48.917 ;
        RECT 43.878 48.889 50.64 48.963 ;
        RECT 43.832 48.935 50.594 49.009 ;
        RECT 43.786 48.981 50.548 49.055 ;
        RECT 43.74 49.027 50.502 49.101 ;
        RECT 43.694 49.073 50.456 49.147 ;
        RECT 43.648 49.119 50.41 49.193 ;
        RECT 43.602 49.165 50.364 49.239 ;
        RECT 43.556 49.211 50.318 49.285 ;
        RECT 43.51 49.257 50.272 49.331 ;
        RECT 43.464 49.303 50.226 49.377 ;
        RECT 43.418 49.349 50.18 49.423 ;
        RECT 43.372 49.395 50.134 49.469 ;
        RECT 43.326 49.441 50.088 49.515 ;
        RECT 43.28 49.487 50.042 49.561 ;
        RECT 43.234 49.533 49.996 49.607 ;
        RECT 43.188 49.579 49.95 49.653 ;
        RECT 43.142 49.625 49.904 49.699 ;
        RECT 43.096 49.671 49.858 49.745 ;
        RECT 43.05 49.717 49.812 49.791 ;
        RECT 43.004 49.763 49.766 49.837 ;
        RECT 42.958 49.809 49.72 49.883 ;
        RECT 42.912 49.855 49.674 49.929 ;
        RECT 42.866 49.901 49.628 49.975 ;
        RECT 42.82 49.947 49.582 50.021 ;
        RECT 42.774 49.993 49.536 50.067 ;
        RECT 42.728 50.039 49.49 50.113 ;
        RECT 42.682 50.085 49.444 50.159 ;
        RECT 42.636 50.131 49.398 50.205 ;
        RECT 42.59 50.177 49.352 50.251 ;
        RECT 42.544 50.223 49.306 50.297 ;
        RECT 42.498 50.269 49.26 50.343 ;
        RECT 42.452 50.315 49.214 50.389 ;
        RECT 42.406 50.361 49.168 50.435 ;
        RECT 42.36 50.407 49.122 50.481 ;
        RECT 42.314 50.453 49.076 50.527 ;
        RECT 42.268 50.499 49.03 50.573 ;
        RECT 42.222 50.545 48.984 50.619 ;
        RECT 42.176 50.591 48.938 50.665 ;
        RECT 42.13 50.637 48.892 50.711 ;
        RECT 42.084 50.683 48.846 50.757 ;
        RECT 42.038 50.729 48.8 50.803 ;
        RECT 41.992 50.775 48.754 50.849 ;
        RECT 41.946 50.821 48.708 50.895 ;
        RECT 41.9 50.867 48.662 50.941 ;
        RECT 41.854 50.913 48.616 50.987 ;
        RECT 41.808 50.959 48.57 51.033 ;
        RECT 41.762 51.005 48.524 51.079 ;
        RECT 41.716 51.051 48.478 51.125 ;
        RECT 41.67 51.097 48.432 51.171 ;
        RECT 41.624 51.143 48.386 51.217 ;
        RECT 41.578 51.189 48.34 51.263 ;
        RECT 41.532 51.235 48.294 51.309 ;
        RECT 41.486 51.281 48.248 51.355 ;
        RECT 41.44 51.327 48.202 51.401 ;
        RECT 41.394 51.373 48.156 51.447 ;
        RECT 41.348 51.419 48.11 51.493 ;
        RECT 41.302 51.465 48.064 51.539 ;
        RECT 41.256 51.511 48.018 51.585 ;
        RECT 41.21 51.557 47.972 51.631 ;
        RECT 41.164 51.603 47.926 51.677 ;
        RECT 41.118 51.649 47.88 51.723 ;
        RECT 41.072 51.695 47.834 51.769 ;
        RECT 41.026 51.741 47.788 51.815 ;
        RECT 40.98 51.787 47.742 51.861 ;
        RECT 40.934 51.833 47.696 51.907 ;
        RECT 40.888 51.879 47.65 51.953 ;
        RECT 40.842 51.925 47.604 51.999 ;
        RECT 40.796 51.971 47.558 52.045 ;
        RECT 40.75 52.017 47.512 52.091 ;
        RECT 40.704 52.063 47.466 52.137 ;
        RECT 40.658 52.109 47.42 52.183 ;
        RECT 40.612 52.155 47.374 52.229 ;
        RECT 40.566 52.201 47.328 52.275 ;
        RECT 40.52 52.247 47.282 52.321 ;
        RECT 40.474 52.293 47.236 52.367 ;
        RECT 40.428 52.339 47.19 52.413 ;
        RECT 40.382 52.385 47.144 52.459 ;
        RECT 40.336 52.431 47.098 52.505 ;
        RECT 40.29 52.477 47.052 52.551 ;
        RECT 40.244 52.523 47.006 52.597 ;
        RECT 40.198 52.569 46.96 52.643 ;
        RECT 40.152 52.615 46.914 52.689 ;
        RECT 40.106 52.661 46.868 52.735 ;
        RECT 40.06 52.707 46.822 52.781 ;
        RECT 40.014 52.753 46.776 52.827 ;
        RECT 39.968 52.799 46.73 52.873 ;
        RECT 39.922 52.845 46.684 52.919 ;
        RECT 39.876 52.891 46.638 52.965 ;
        RECT 39.83 52.937 46.592 53.011 ;
        RECT 39.784 52.983 46.546 53.057 ;
        RECT 39.738 53.029 46.5 53.103 ;
        RECT 39.692 53.075 46.454 53.149 ;
        RECT 39.646 53.121 46.408 53.195 ;
        RECT 39.6 53.167 46.362 53.241 ;
        RECT 39.554 53.213 46.316 53.287 ;
        RECT 39.508 53.259 46.27 53.333 ;
        RECT 39.462 53.305 46.224 53.379 ;
        RECT 39.416 53.351 46.178 53.425 ;
        RECT 39.37 53.397 46.132 53.471 ;
        RECT 39.324 53.443 46.086 53.517 ;
        RECT 39.278 53.489 46.04 53.563 ;
        RECT 39.232 53.535 45.994 53.609 ;
        RECT 39.186 53.581 45.948 53.655 ;
        RECT 39.14 53.627 45.902 53.701 ;
        RECT 39.094 53.673 45.856 53.747 ;
        RECT 39.048 53.719 45.81 53.793 ;
        RECT 39.002 53.765 45.764 53.839 ;
        RECT 38.956 53.811 45.718 53.885 ;
        RECT 38.91 53.857 45.672 53.931 ;
        RECT 38.864 53.903 45.626 53.977 ;
        RECT 38.818 53.949 45.58 54.023 ;
        RECT 38.772 53.995 45.534 54.069 ;
        RECT 38.726 54.041 45.488 54.115 ;
        RECT 38.68 54.087 45.442 54.161 ;
        RECT 38.634 54.133 45.396 54.207 ;
        RECT 38.588 54.179 45.35 54.253 ;
        RECT 38.542 54.225 45.304 54.299 ;
        RECT 38.496 54.271 45.258 54.345 ;
        RECT 38.45 54.317 45.212 54.391 ;
        RECT 38.404 54.363 45.166 54.437 ;
        RECT 38.358 54.409 45.12 54.483 ;
        RECT 38.312 54.455 45.074 54.529 ;
        RECT 38.266 54.501 45.028 54.575 ;
        RECT 38.22 54.547 44.982 54.621 ;
        RECT 38.174 54.593 44.936 54.667 ;
        RECT 38.128 54.639 44.89 54.713 ;
        RECT 38.082 54.685 44.844 54.759 ;
        RECT 38.036 54.731 44.798 54.805 ;
        RECT 37.99 54.777 44.752 54.851 ;
        RECT 37.944 54.823 44.706 54.897 ;
        RECT 37.898 54.869 44.66 54.943 ;
        RECT 37.852 54.915 44.614 54.989 ;
        RECT 37.806 54.961 44.568 55.035 ;
        RECT 37.76 55.007 44.522 55.081 ;
        RECT 37.714 55.053 44.476 55.127 ;
        RECT 37.668 55.099 44.43 55.173 ;
        RECT 37.622 55.145 44.384 55.219 ;
        RECT 37.576 55.191 44.338 55.265 ;
        RECT 37.53 55.237 44.292 55.311 ;
        RECT 37.484 55.283 44.246 55.357 ;
        RECT 37.438 55.329 44.2 55.403 ;
        RECT 37.392 55.375 44.154 55.449 ;
        RECT 37.346 55.421 44.108 55.495 ;
        RECT 37.3 55.467 44.062 55.541 ;
        RECT 37.254 55.513 44.016 55.587 ;
        RECT 37.208 55.559 43.97 55.633 ;
        RECT 37.162 55.605 43.924 55.679 ;
        RECT 37.116 55.651 43.878 55.725 ;
        RECT 37.07 55.697 43.832 55.771 ;
        RECT 37.024 55.743 43.786 55.817 ;
        RECT 36.978 55.789 43.74 55.863 ;
        RECT 36.932 55.835 43.694 55.909 ;
        RECT 36.886 55.881 43.648 55.955 ;
        RECT 36.84 55.927 43.602 56.001 ;
        RECT 36.794 55.973 43.556 56.047 ;
        RECT 36.748 56.019 43.51 56.093 ;
        RECT 36.702 56.065 43.464 56.139 ;
        RECT 36.656 56.111 43.418 56.185 ;
        RECT 36.61 56.157 43.372 56.231 ;
        RECT 36.564 56.203 43.326 56.277 ;
        RECT 36.518 56.249 43.28 56.323 ;
        RECT 36.472 56.295 43.234 56.369 ;
        RECT 36.426 56.341 43.188 56.415 ;
        RECT 36.38 56.387 43.142 56.461 ;
        RECT 36.334 56.433 43.096 56.507 ;
        RECT 36.288 56.479 43.05 56.553 ;
        RECT 36.242 56.525 43.004 56.599 ;
        RECT 36.196 56.571 42.958 56.645 ;
        RECT 36.15 56.617 42.912 56.691 ;
        RECT 36.104 56.663 42.866 56.737 ;
        RECT 36.058 56.709 42.82 56.783 ;
        RECT 36.012 56.755 42.774 56.829 ;
        RECT 35.966 56.801 42.728 56.875 ;
        RECT 35.92 56.847 42.682 56.921 ;
        RECT 35.874 56.893 42.636 56.967 ;
        RECT 35.828 56.939 42.59 57.013 ;
        RECT 35.782 56.985 42.544 57.059 ;
        RECT 35.736 57.031 42.498 57.105 ;
        RECT 35.69 57.077 42.452 57.151 ;
        RECT 35.644 57.123 42.406 57.197 ;
        RECT 35.598 57.169 42.36 57.243 ;
        RECT 35.552 57.215 42.314 57.289 ;
        RECT 35.506 57.261 42.268 57.335 ;
        RECT 35.46 57.307 42.222 57.381 ;
        RECT 35.414 57.353 42.176 57.427 ;
        RECT 35.368 57.399 42.13 57.473 ;
        RECT 35.322 57.445 42.084 57.519 ;
        RECT 35.276 57.491 42.038 57.565 ;
        RECT 35.23 57.537 41.992 57.611 ;
        RECT 35.184 57.583 41.946 57.657 ;
        RECT 35.138 57.629 41.9 57.703 ;
        RECT 35.092 57.675 41.854 57.749 ;
        RECT 35.046 57.721 41.808 57.795 ;
        RECT 34.984 57.798 41.762 57.841 ;
        RECT 35 57.767 41.762 57.841 ;
        RECT 34.938 57.829 41.716 57.887 ;
        RECT 34.892 57.875 41.67 57.933 ;
        RECT 34.846 57.921 41.624 57.979 ;
        RECT 34.8 57.967 41.578 58.025 ;
        RECT 34.754 58.013 41.532 58.071 ;
        RECT 34.708 58.059 41.486 58.117 ;
        RECT 34.662 58.105 41.44 58.163 ;
        RECT 34.616 58.151 41.394 58.209 ;
        RECT 34.57 58.197 41.348 58.255 ;
        RECT 34.524 58.243 41.302 58.301 ;
        RECT 34.478 58.289 41.256 58.347 ;
        RECT 34.432 58.335 41.21 58.393 ;
        RECT 34.386 58.381 41.164 58.439 ;
        RECT 34.34 58.427 41.118 58.485 ;
        RECT 34.294 58.473 41.072 58.531 ;
        RECT 34.248 58.519 41.026 58.577 ;
        RECT 34.202 58.565 40.98 58.623 ;
        RECT 34.156 58.611 40.934 58.669 ;
        RECT 34.11 58.657 40.888 58.715 ;
        RECT 34.064 58.703 40.842 58.761 ;
        RECT 34.018 58.749 40.796 58.807 ;
        RECT 33.972 58.795 40.75 58.853 ;
        RECT 33.926 58.841 40.704 58.899 ;
        RECT 33.88 58.887 40.658 58.945 ;
        RECT 33.834 58.933 40.612 58.991 ;
        RECT 33.788 58.979 40.566 59.037 ;
        RECT 33.742 59.025 40.52 59.083 ;
        RECT 33.696 59.071 40.474 59.129 ;
        RECT 33.65 59.117 40.428 59.175 ;
        RECT 33.604 59.163 40.382 59.221 ;
        RECT 33.558 59.209 40.336 59.267 ;
        RECT 33.512 59.255 40.29 59.313 ;
        RECT 33.466 59.301 40.244 59.359 ;
        RECT 33.42 59.347 40.198 59.405 ;
        RECT 33.374 59.393 40.152 59.451 ;
        RECT 33.328 59.439 40.106 59.497 ;
        RECT 33.282 59.485 40.06 59.543 ;
        RECT 33.236 59.531 40.014 59.589 ;
        RECT 33.19 59.577 39.968 59.635 ;
        RECT 33.144 59.623 39.922 59.681 ;
        RECT 33.098 59.669 39.876 59.727 ;
        RECT 33.052 59.715 39.83 59.773 ;
        RECT 33.006 59.761 39.784 59.819 ;
        RECT 32.96 59.807 39.738 59.865 ;
        RECT 32.914 59.853 39.692 59.911 ;
        RECT 32.868 59.899 39.646 59.957 ;
        RECT 32.822 59.945 39.6 60.003 ;
        RECT 32.776 59.991 39.554 60.049 ;
        RECT 32.73 60.037 39.508 60.095 ;
        RECT 32.684 60.083 39.462 60.141 ;
        RECT 32.638 60.129 39.416 60.187 ;
        RECT 32.592 60.175 39.37 60.233 ;
        RECT 32.546 60.221 39.324 60.279 ;
        RECT 32.5 60.267 39.278 60.325 ;
        RECT 32.454 60.313 39.232 60.371 ;
        RECT 32.408 60.359 39.186 60.417 ;
        RECT 32.362 60.405 39.14 60.463 ;
        RECT 32.316 60.451 39.094 60.509 ;
        RECT 32.27 60.497 39.048 60.555 ;
        RECT 32.224 60.543 39.002 60.601 ;
        RECT 32.178 60.589 38.956 60.647 ;
        RECT 32.132 60.635 38.91 60.693 ;
        RECT 32.086 60.681 38.864 60.739 ;
        RECT 32.04 60.727 38.818 60.785 ;
        RECT 31.994 60.773 38.772 60.831 ;
        RECT 31.948 60.819 38.726 60.877 ;
        RECT 31.902 60.865 38.68 60.923 ;
        RECT 31.856 60.911 38.634 60.969 ;
        RECT 31.81 60.957 38.588 61.015 ;
        RECT 31.764 61.003 38.542 61.061 ;
        RECT 31.718 61.049 38.496 61.107 ;
        RECT 31.672 61.095 38.45 61.153 ;
        RECT 31.626 61.141 38.404 61.199 ;
        RECT 31.58 61.187 38.358 61.245 ;
        RECT 31.534 61.233 38.312 61.291 ;
        RECT 31.488 61.279 38.266 61.337 ;
        RECT 31.442 61.325 38.22 61.383 ;
        RECT 31.396 61.371 38.174 61.429 ;
        RECT 31.35 61.417 38.128 61.475 ;
        RECT 31.304 61.463 38.082 61.521 ;
        RECT 31.258 61.509 38.036 61.567 ;
        RECT 31.212 61.555 37.99 61.613 ;
        RECT 31.166 61.601 37.944 61.659 ;
        RECT 31.12 61.647 37.898 61.705 ;
        RECT 31.074 61.693 37.852 61.751 ;
        RECT 31.028 61.739 37.806 61.797 ;
        RECT 30.982 61.785 37.76 61.843 ;
        RECT 30.936 61.831 37.714 61.889 ;
        RECT 30.89 61.877 37.668 61.935 ;
        RECT 30.844 61.923 37.622 61.981 ;
        RECT 30.798 61.969 37.576 62.027 ;
        RECT 30.752 62.015 37.53 62.073 ;
        RECT 30.706 62.061 37.484 62.119 ;
        RECT 30.66 62.107 37.438 62.165 ;
        RECT 30.614 62.153 37.392 62.211 ;
        RECT 30.568 62.199 37.346 62.257 ;
        RECT 30.522 62.245 37.3 62.303 ;
        RECT 30.476 62.291 37.254 62.349 ;
        RECT 30.43 62.337 37.208 62.395 ;
        RECT 30.384 62.383 37.162 62.441 ;
        RECT 30.338 62.429 37.116 62.487 ;
        RECT 30.292 62.475 37.07 62.533 ;
        RECT 30.246 62.521 37.024 62.579 ;
        RECT 30.2 62.567 36.978 62.625 ;
        RECT 30.2 62.567 36.932 62.671 ;
        RECT 30.2 62.567 36.886 62.717 ;
        RECT 30.2 62.567 36.84 62.763 ;
        RECT 30.2 62.567 36.794 62.809 ;
        RECT 30.2 62.567 36.748 62.855 ;
        RECT 30.2 62.567 36.702 62.901 ;
        RECT 30.2 62.567 36.656 62.947 ;
        RECT 30.2 62.567 36.61 62.993 ;
        RECT 30.2 62.567 36.564 63.039 ;
        RECT 30.2 62.567 36.518 63.085 ;
        RECT 30.2 62.567 36.472 63.131 ;
        RECT 30.2 62.567 36.426 63.177 ;
        RECT 30.2 62.567 36.38 63.223 ;
        RECT 30.2 62.567 36.334 63.269 ;
        RECT 30.2 62.567 36.288 63.315 ;
        RECT 30.2 62.567 36.242 63.361 ;
        RECT 30.2 62.567 36.196 63.407 ;
        RECT 30.2 62.567 36.15 63.453 ;
        RECT 30.2 62.567 36.104 63.499 ;
        RECT 30.2 62.567 36.058 63.545 ;
        RECT 30.2 62.567 36.012 63.591 ;
        RECT 30.2 62.567 35.966 63.637 ;
        RECT 30.2 62.567 35.92 63.683 ;
        RECT 30.2 62.567 35.874 63.729 ;
        RECT 30.2 62.567 35.828 63.775 ;
        RECT 30.2 62.567 35.782 63.821 ;
        RECT 30.2 62.567 35.736 63.867 ;
        RECT 30.2 62.567 35.69 63.913 ;
        RECT 30.2 62.567 35.644 63.959 ;
        RECT 30.2 62.567 35.598 64.005 ;
        RECT 30.2 62.567 35.552 64.051 ;
        RECT 30.2 62.567 35.506 64.097 ;
        RECT 30.2 62.567 35.46 64.143 ;
        RECT 30.2 62.567 35.414 64.189 ;
        RECT 30.2 62.567 35.368 64.235 ;
        RECT 30.2 62.567 35.322 64.281 ;
        RECT 30.2 62.567 35.276 64.327 ;
        RECT 30.2 62.567 35.23 64.373 ;
        RECT 30.2 62.567 35.184 64.419 ;
        RECT 30.2 62.567 35.138 64.465 ;
        RECT 30.2 62.567 35.092 64.511 ;
        RECT 30.2 62.567 35.046 64.557 ;
        RECT 30.2 62.567 35 80 ;
    END
    PORT
      LAYER QB ;
        RECT 17.734 57.493 24.496 57.567 ;
        RECT 17.688 57.539 24.45 57.613 ;
        RECT 17.642 57.585 24.404 57.659 ;
        RECT 17.596 57.631 24.358 57.705 ;
        RECT 17.55 57.677 24.312 57.751 ;
        RECT 17.504 57.723 24.266 57.797 ;
        RECT 17.458 57.769 24.22 57.843 ;
        RECT 17.412 57.815 24.174 57.889 ;
        RECT 17.366 57.861 24.128 57.935 ;
        RECT 17.32 57.907 24.082 57.981 ;
        RECT 17.274 57.953 24.036 58.027 ;
        RECT 17.228 57.999 23.99 58.073 ;
        RECT 17.182 58.045 23.944 58.119 ;
        RECT 17.136 58.091 23.898 58.165 ;
        RECT 17.09 58.137 23.852 58.211 ;
        RECT 17.044 58.183 23.806 58.257 ;
        RECT 16.998 58.229 23.76 58.303 ;
        RECT 16.952 58.275 23.714 58.349 ;
        RECT 16.906 58.321 23.668 58.395 ;
        RECT 16.86 58.367 23.622 58.441 ;
        RECT 16.814 58.413 23.576 58.487 ;
        RECT 16.768 58.459 23.53 58.533 ;
        RECT 16.722 58.505 23.484 58.579 ;
        RECT 16.676 58.551 23.438 58.625 ;
        RECT 16.63 58.597 23.392 58.671 ;
        RECT 16.584 58.643 23.346 58.717 ;
        RECT 16.538 58.689 23.3 58.763 ;
        RECT 16.492 58.735 23.254 58.809 ;
        RECT 16.446 58.781 23.208 58.855 ;
        RECT 16.384 58.858 23.162 58.901 ;
        RECT 16.4 58.827 23.162 58.901 ;
        RECT 16.338 58.889 23.116 58.947 ;
        RECT 16.292 58.935 23.07 58.993 ;
        RECT 16.246 58.981 23.024 59.039 ;
        RECT 16.2 59.027 22.978 59.085 ;
        RECT 16.154 59.073 22.932 59.131 ;
        RECT 16.108 59.119 22.886 59.177 ;
        RECT 16.062 59.165 22.84 59.223 ;
        RECT 16.016 59.211 22.794 59.269 ;
        RECT 15.97 59.257 22.748 59.315 ;
        RECT 15.924 59.303 22.702 59.361 ;
        RECT 15.878 59.349 22.656 59.407 ;
        RECT 15.832 59.395 22.61 59.453 ;
        RECT 15.786 59.441 22.564 59.499 ;
        RECT 15.74 59.487 22.518 59.545 ;
        RECT 15.694 59.533 22.472 59.591 ;
        RECT 15.648 59.579 22.426 59.637 ;
        RECT 15.602 59.625 22.38 59.683 ;
        RECT 15.556 59.671 22.334 59.729 ;
        RECT 15.51 59.717 22.288 59.775 ;
        RECT 15.464 59.763 22.242 59.821 ;
        RECT 15.418 59.809 22.196 59.867 ;
        RECT 15.372 59.855 22.15 59.913 ;
        RECT 15.326 59.901 22.104 59.959 ;
        RECT 15.28 59.947 22.058 60.005 ;
        RECT 15.234 59.993 22.012 60.051 ;
        RECT 15.188 60.039 21.966 60.097 ;
        RECT 15.142 60.085 21.92 60.143 ;
        RECT 15.096 60.131 21.874 60.189 ;
        RECT 15.05 60.177 21.828 60.235 ;
        RECT 15.004 60.223 21.782 60.281 ;
        RECT 14.958 60.269 21.736 60.327 ;
        RECT 14.912 60.315 21.69 60.373 ;
        RECT 14.866 60.361 21.644 60.419 ;
        RECT 14.82 60.407 21.598 60.465 ;
        RECT 14.774 60.453 21.552 60.511 ;
        RECT 14.728 60.499 21.506 60.557 ;
        RECT 14.682 60.545 21.46 60.603 ;
        RECT 14.636 60.591 21.414 60.649 ;
        RECT 14.59 60.637 21.368 60.695 ;
        RECT 14.544 60.683 21.322 60.741 ;
        RECT 14.498 60.729 21.276 60.787 ;
        RECT 14.452 60.775 21.23 60.833 ;
        RECT 14.406 60.821 21.184 60.879 ;
        RECT 14.36 60.867 21.138 60.925 ;
        RECT 14.314 60.913 21.092 60.971 ;
        RECT 14.268 60.959 21.046 61.017 ;
        RECT 14.222 61.005 21 61.063 ;
        RECT 14.176 61.051 20.954 61.109 ;
        RECT 14.13 61.097 20.908 61.155 ;
        RECT 14.084 61.143 20.862 61.201 ;
        RECT 14.038 61.189 20.816 61.247 ;
        RECT 13.992 61.235 20.77 61.293 ;
        RECT 13.946 61.281 20.724 61.339 ;
        RECT 13.9 61.327 20.678 61.385 ;
        RECT 13.854 61.373 20.632 61.431 ;
        RECT 13.808 61.419 20.586 61.477 ;
        RECT 13.762 61.465 20.54 61.523 ;
        RECT 13.716 61.511 20.494 61.569 ;
        RECT 13.67 61.557 20.448 61.615 ;
        RECT 13.624 61.603 20.402 61.661 ;
        RECT 13.578 61.649 20.356 61.707 ;
        RECT 13.532 61.695 20.31 61.753 ;
        RECT 13.486 61.741 20.264 61.799 ;
        RECT 13.44 61.787 20.218 61.845 ;
        RECT 13.394 61.833 20.172 61.891 ;
        RECT 13.348 61.879 20.126 61.937 ;
        RECT 13.302 61.925 20.08 61.983 ;
        RECT 13.256 61.971 20.034 62.029 ;
        RECT 13.21 62.017 19.988 62.075 ;
        RECT 13.164 62.063 19.942 62.121 ;
        RECT 13.118 62.109 19.896 62.167 ;
        RECT 13.072 62.155 19.85 62.213 ;
        RECT 13.026 62.201 19.804 62.259 ;
        RECT 12.98 62.247 19.758 62.305 ;
        RECT 12.934 62.293 19.712 62.351 ;
        RECT 12.888 62.339 19.666 62.397 ;
        RECT 12.842 62.385 19.62 62.443 ;
        RECT 12.796 62.431 19.574 62.489 ;
        RECT 12.75 62.477 19.528 62.535 ;
        RECT 12.704 62.523 19.482 62.581 ;
        RECT 12.658 62.569 19.436 62.627 ;
        RECT 12.612 62.615 19.39 62.673 ;
        RECT 12.566 62.661 19.344 62.719 ;
        RECT 12.52 62.707 19.298 62.765 ;
        RECT 12.474 62.753 19.252 62.811 ;
        RECT 12.428 62.799 19.206 62.857 ;
        RECT 12.382 62.845 19.16 62.903 ;
        RECT 12.336 62.891 19.114 62.949 ;
        RECT 12.29 62.937 19.068 62.995 ;
        RECT 12.244 62.983 19.022 63.041 ;
        RECT 12.198 63.029 18.976 63.087 ;
        RECT 12.152 63.075 18.93 63.133 ;
        RECT 12.106 63.121 18.884 63.179 ;
        RECT 12.06 63.167 18.838 63.225 ;
        RECT 12.014 63.213 18.792 63.271 ;
        RECT 11.968 63.259 18.746 63.317 ;
        RECT 11.922 63.305 18.7 63.363 ;
        RECT 11.876 63.351 18.654 63.409 ;
        RECT 11.83 63.397 18.608 63.455 ;
        RECT 11.784 63.443 18.562 63.501 ;
        RECT 11.738 63.489 18.516 63.547 ;
        RECT 11.692 63.535 18.47 63.593 ;
        RECT 11.646 63.581 18.424 63.639 ;
        RECT 11.6 63.627 18.378 63.685 ;
        RECT 11.6 63.627 18.332 63.731 ;
        RECT 11.6 63.627 18.286 63.777 ;
        RECT 11.6 63.627 18.24 63.823 ;
        RECT 11.6 63.627 18.194 63.869 ;
        RECT 11.6 63.627 18.148 63.915 ;
        RECT 11.6 63.627 18.102 63.961 ;
        RECT 11.6 63.627 18.056 64.007 ;
        RECT 11.6 63.627 18.01 64.053 ;
        RECT 11.6 63.627 17.964 64.099 ;
        RECT 11.6 63.627 17.918 64.145 ;
        RECT 11.6 63.627 17.872 64.191 ;
        RECT 11.6 63.627 17.826 64.237 ;
        RECT 11.6 63.627 17.78 64.283 ;
        RECT 11.6 63.627 17.734 64.329 ;
        RECT 11.6 63.627 17.688 64.375 ;
        RECT 11.6 63.627 17.642 64.421 ;
        RECT 11.6 63.627 17.596 64.467 ;
        RECT 11.6 63.627 17.55 64.513 ;
        RECT 11.6 63.627 17.504 64.559 ;
        RECT 11.6 63.627 17.458 64.605 ;
        RECT 11.6 63.627 17.412 64.651 ;
        RECT 11.6 63.627 17.366 64.697 ;
        RECT 11.6 63.627 17.32 64.743 ;
        RECT 11.6 63.627 17.274 64.789 ;
        RECT 11.6 63.627 17.228 64.835 ;
        RECT 11.6 63.627 17.182 64.881 ;
        RECT 11.6 63.627 17.136 64.927 ;
        RECT 11.6 63.627 17.09 64.973 ;
        RECT 11.6 63.627 17.044 65.019 ;
        RECT 11.6 63.627 16.998 65.065 ;
        RECT 11.6 63.627 16.952 65.111 ;
        RECT 11.6 63.627 16.906 65.157 ;
        RECT 11.6 63.627 16.86 65.203 ;
        RECT 11.6 63.627 16.814 65.249 ;
        RECT 11.6 63.627 16.768 65.295 ;
        RECT 11.6 63.627 16.722 65.341 ;
        RECT 11.6 63.627 16.676 65.387 ;
        RECT 11.6 63.627 16.63 65.433 ;
        RECT 11.6 63.627 16.584 65.479 ;
        RECT 11.6 63.627 16.538 65.525 ;
        RECT 11.6 63.627 16.492 65.571 ;
        RECT 11.6 63.627 16.446 65.617 ;
        RECT 11.6 63.627 16.4 80 ;
        RECT 63.65 11.6 80 16.4 ;
        RECT 58.858 16.369 65.64 16.406 ;
        RECT 56.88 18.347 63.65 18.394 ;
        RECT 56.926 18.301 63.696 18.367 ;
        RECT 63.642 11.604 63.65 18.394 ;
        RECT 56.972 18.255 63.742 18.321 ;
        RECT 63.596 11.631 63.642 18.421 ;
        RECT 56.834 18.393 63.596 18.467 ;
        RECT 57.018 18.209 63.788 18.275 ;
        RECT 63.55 11.677 63.596 18.467 ;
        RECT 56.788 18.439 63.55 18.513 ;
        RECT 57.064 18.163 63.834 18.229 ;
        RECT 63.504 11.723 63.55 18.513 ;
        RECT 56.742 18.485 63.504 18.559 ;
        RECT 57.11 18.117 63.88 18.183 ;
        RECT 63.458 11.769 63.504 18.559 ;
        RECT 56.696 18.531 63.458 18.605 ;
        RECT 57.156 18.071 63.926 18.137 ;
        RECT 63.412 11.815 63.458 18.605 ;
        RECT 56.65 18.577 63.412 18.651 ;
        RECT 57.202 18.025 63.972 18.091 ;
        RECT 63.366 11.861 63.412 18.651 ;
        RECT 56.604 18.623 63.366 18.697 ;
        RECT 57.248 17.979 64.018 18.045 ;
        RECT 63.32 11.907 63.366 18.697 ;
        RECT 56.558 18.669 63.32 18.743 ;
        RECT 57.294 17.933 64.064 17.999 ;
        RECT 63.274 11.953 63.32 18.743 ;
        RECT 56.512 18.715 63.274 18.789 ;
        RECT 57.34 17.887 64.11 17.953 ;
        RECT 63.228 11.999 63.274 18.789 ;
        RECT 56.466 18.761 63.228 18.835 ;
        RECT 57.386 17.841 64.156 17.907 ;
        RECT 63.182 12.045 63.228 18.835 ;
        RECT 56.42 18.807 63.182 18.881 ;
        RECT 57.432 17.795 64.202 17.861 ;
        RECT 63.136 12.091 63.182 18.881 ;
        RECT 56.374 18.853 63.136 18.927 ;
        RECT 57.478 17.749 64.248 17.815 ;
        RECT 63.09 12.137 63.136 18.927 ;
        RECT 56.328 18.899 63.09 18.973 ;
        RECT 57.524 17.703 64.294 17.769 ;
        RECT 63.044 12.183 63.09 18.973 ;
        RECT 56.282 18.945 63.044 19.019 ;
        RECT 57.57 17.657 64.34 17.723 ;
        RECT 62.998 12.229 63.044 19.019 ;
        RECT 56.236 18.991 62.998 19.065 ;
        RECT 57.616 17.611 64.386 17.677 ;
        RECT 62.952 12.275 62.998 19.065 ;
        RECT 56.19 19.037 62.952 19.111 ;
        RECT 57.662 17.565 64.432 17.631 ;
        RECT 62.906 12.321 62.952 19.111 ;
        RECT 56.144 19.083 62.906 19.157 ;
        RECT 57.708 17.519 64.478 17.585 ;
        RECT 62.86 12.367 62.906 19.157 ;
        RECT 56.098 19.129 62.86 19.203 ;
        RECT 57.754 17.473 64.524 17.539 ;
        RECT 62.814 12.413 62.86 19.203 ;
        RECT 56.052 19.175 62.814 19.249 ;
        RECT 57.8 17.427 64.57 17.493 ;
        RECT 62.768 12.459 62.814 19.249 ;
        RECT 56.006 19.221 62.768 19.295 ;
        RECT 57.846 17.381 64.616 17.447 ;
        RECT 62.722 12.505 62.768 19.295 ;
        RECT 55.96 19.267 62.722 19.341 ;
        RECT 57.892 17.335 64.662 17.401 ;
        RECT 62.676 12.551 62.722 19.341 ;
        RECT 55.914 19.313 62.676 19.387 ;
        RECT 57.938 17.289 64.708 17.355 ;
        RECT 62.63 12.597 62.676 19.387 ;
        RECT 55.868 19.359 62.63 19.433 ;
        RECT 57.984 17.243 64.754 17.309 ;
        RECT 62.584 12.643 62.63 19.433 ;
        RECT 55.822 19.405 62.584 19.479 ;
        RECT 58.03 17.197 64.8 17.263 ;
        RECT 62.538 12.689 62.584 19.479 ;
        RECT 55.776 19.451 62.538 19.525 ;
        RECT 58.076 17.151 64.846 17.217 ;
        RECT 62.492 12.735 62.538 19.525 ;
        RECT 55.73 19.497 62.492 19.571 ;
        RECT 58.122 17.105 64.892 17.171 ;
        RECT 62.446 12.781 62.492 19.571 ;
        RECT 55.684 19.543 62.446 19.617 ;
        RECT 58.168 17.059 64.938 17.125 ;
        RECT 62.4 12.827 62.446 19.617 ;
        RECT 55.638 19.589 62.4 19.663 ;
        RECT 58.214 17.013 64.984 17.079 ;
        RECT 62.354 12.873 62.4 19.663 ;
        RECT 55.592 19.635 62.354 19.709 ;
        RECT 58.26 16.967 65.03 17.033 ;
        RECT 62.308 12.919 62.354 19.709 ;
        RECT 55.546 19.681 62.308 19.755 ;
        RECT 58.306 16.921 65.076 16.987 ;
        RECT 62.262 12.965 62.308 19.755 ;
        RECT 55.5 19.727 62.262 19.801 ;
        RECT 58.352 16.875 65.122 16.941 ;
        RECT 62.216 13.011 62.262 19.801 ;
        RECT 55.454 19.773 62.216 19.847 ;
        RECT 58.398 16.829 65.168 16.895 ;
        RECT 62.17 13.057 62.216 19.847 ;
        RECT 55.408 19.819 62.17 19.893 ;
        RECT 58.444 16.783 65.214 16.849 ;
        RECT 62.124 13.103 62.17 19.893 ;
        RECT 55.362 19.865 62.124 19.939 ;
        RECT 58.49 16.737 65.26 16.803 ;
        RECT 62.078 13.149 62.124 19.939 ;
        RECT 55.316 19.911 62.078 19.985 ;
        RECT 58.536 16.691 65.306 16.757 ;
        RECT 62.032 13.195 62.078 19.985 ;
        RECT 55.27 19.957 62.032 20.031 ;
        RECT 58.582 16.645 65.352 16.711 ;
        RECT 61.986 13.241 62.032 20.031 ;
        RECT 55.224 20.003 61.986 20.077 ;
        RECT 58.628 16.599 65.398 16.665 ;
        RECT 61.94 13.287 61.986 20.077 ;
        RECT 55.178 20.049 61.94 20.123 ;
        RECT 58.674 16.553 65.444 16.619 ;
        RECT 61.894 13.333 61.94 20.123 ;
        RECT 55.132 20.095 61.894 20.169 ;
        RECT 58.72 16.507 65.49 16.573 ;
        RECT 61.848 13.379 61.894 20.169 ;
        RECT 55.086 20.141 61.848 20.215 ;
        RECT 58.766 16.461 65.536 16.527 ;
        RECT 61.802 13.425 61.848 20.215 ;
        RECT 55.04 20.187 61.802 20.261 ;
        RECT 58.812 16.415 65.582 16.481 ;
        RECT 61.756 13.471 61.802 20.261 ;
        RECT 54.994 20.233 61.756 20.307 ;
        RECT 58.858 16.369 65.628 16.435 ;
        RECT 61.71 13.517 61.756 20.307 ;
        RECT 54.948 20.279 61.71 20.353 ;
        RECT 58.904 16.323 80 16.4 ;
        RECT 61.664 13.563 61.71 20.353 ;
        RECT 54.902 20.325 61.664 20.399 ;
        RECT 58.95 16.277 80 16.4 ;
        RECT 61.618 13.609 61.664 20.399 ;
        RECT 54.856 20.371 61.618 20.445 ;
        RECT 58.996 16.231 80 16.4 ;
        RECT 61.572 13.655 61.618 20.445 ;
        RECT 54.81 20.417 61.572 20.491 ;
        RECT 59.042 16.185 80 16.4 ;
        RECT 61.526 13.701 61.572 20.491 ;
        RECT 54.764 20.463 61.526 20.537 ;
        RECT 59.088 16.139 80 16.4 ;
        RECT 61.48 13.747 61.526 20.537 ;
        RECT 54.718 20.509 61.48 20.583 ;
        RECT 59.134 16.093 80 16.4 ;
        RECT 61.434 13.793 61.48 20.583 ;
        RECT 54.672 20.555 61.434 20.629 ;
        RECT 59.18 16.047 80 16.4 ;
        RECT 61.388 13.839 61.434 20.629 ;
        RECT 54.626 20.601 61.388 20.675 ;
        RECT 59.226 16.001 80 16.4 ;
        RECT 61.342 13.885 61.388 20.675 ;
        RECT 54.58 20.647 61.342 20.721 ;
        RECT 59.272 15.955 80 16.4 ;
        RECT 61.296 13.931 61.342 20.721 ;
        RECT 54.534 20.693 61.296 20.767 ;
        RECT 59.318 15.909 80 16.4 ;
        RECT 61.25 13.977 61.296 20.767 ;
        RECT 54.488 20.739 61.25 20.813 ;
        RECT 59.364 15.863 80 16.4 ;
        RECT 61.204 14.023 61.25 20.813 ;
        RECT 54.442 20.785 61.204 20.859 ;
        RECT 59.41 15.817 80 16.4 ;
        RECT 61.158 14.069 61.204 20.859 ;
        RECT 54.396 20.831 61.158 20.905 ;
        RECT 59.456 15.771 80 16.4 ;
        RECT 61.112 14.115 61.158 20.905 ;
        RECT 54.35 20.877 61.112 20.951 ;
        RECT 59.502 15.725 80 16.4 ;
        RECT 61.066 14.161 61.112 20.951 ;
        RECT 54.304 20.923 61.066 20.997 ;
        RECT 59.548 15.679 80 16.4 ;
        RECT 61.02 14.207 61.066 20.997 ;
        RECT 54.258 20.969 61.02 21.043 ;
        RECT 59.594 15.633 80 16.4 ;
        RECT 60.974 14.253 61.02 21.043 ;
        RECT 54.212 21.015 60.974 21.089 ;
        RECT 59.64 15.587 80 16.4 ;
        RECT 60.928 14.299 60.974 21.089 ;
        RECT 54.166 21.061 60.928 21.135 ;
        RECT 59.686 15.541 80 16.4 ;
        RECT 60.882 14.345 60.928 21.135 ;
        RECT 54.12 21.107 60.882 21.181 ;
        RECT 59.732 15.495 80 16.4 ;
        RECT 60.836 14.391 60.882 21.181 ;
        RECT 54.074 21.153 60.836 21.227 ;
        RECT 59.778 15.449 80 16.4 ;
        RECT 60.79 14.437 60.836 21.227 ;
        RECT 54.028 21.199 60.79 21.273 ;
        RECT 59.824 15.403 80 16.4 ;
        RECT 60.744 14.483 60.79 21.273 ;
        RECT 53.982 21.245 60.744 21.319 ;
        RECT 59.87 15.357 80 16.4 ;
        RECT 60.698 14.529 60.744 21.319 ;
        RECT 53.936 21.291 60.698 21.365 ;
        RECT 59.916 15.311 80 16.4 ;
        RECT 60.652 14.575 60.698 21.365 ;
        RECT 53.89 21.337 60.652 21.411 ;
        RECT 59.962 15.265 80 16.4 ;
        RECT 60.606 14.621 60.652 21.411 ;
        RECT 53.844 21.383 60.606 21.457 ;
        RECT 60.008 15.219 80 16.4 ;
        RECT 60.56 14.667 60.606 21.457 ;
        RECT 53.798 21.429 60.56 21.503 ;
        RECT 60.054 15.173 80 16.4 ;
        RECT 60.514 14.713 60.56 21.503 ;
        RECT 53.752 21.475 60.514 21.549 ;
        RECT 60.1 15.127 80 16.4 ;
        RECT 60.468 14.759 60.514 21.549 ;
        RECT 53.706 21.521 60.468 21.595 ;
        RECT 60.146 15.081 80 16.4 ;
        RECT 60.422 14.805 60.468 21.595 ;
        RECT 53.66 21.567 60.422 21.641 ;
        RECT 60.192 15.035 80 16.4 ;
        RECT 60.376 14.851 60.422 21.641 ;
        RECT 53.614 21.613 60.376 21.687 ;
        RECT 60.238 14.989 80 16.4 ;
        RECT 60.33 14.897 60.376 21.687 ;
        RECT 53.568 21.659 60.33 21.733 ;
        RECT 60.284 14.943 80 16.4 ;
        RECT 53.522 21.705 60.284 21.779 ;
        RECT 53.476 21.751 60.238 21.825 ;
        RECT 53.43 21.797 60.192 21.871 ;
        RECT 53.384 21.843 60.146 21.917 ;
        RECT 53.338 21.889 60.1 21.963 ;
        RECT 53.292 21.935 60.054 22.009 ;
        RECT 53.246 21.981 60.008 22.055 ;
        RECT 53.2 22.027 59.962 22.101 ;
        RECT 53.154 22.073 59.916 22.147 ;
        RECT 53.108 22.119 59.87 22.193 ;
        RECT 53.062 22.165 59.824 22.239 ;
        RECT 53.016 22.211 59.778 22.285 ;
        RECT 52.97 22.257 59.732 22.331 ;
        RECT 52.924 22.303 59.686 22.377 ;
        RECT 52.878 22.349 59.64 22.423 ;
        RECT 52.832 22.395 59.594 22.469 ;
        RECT 52.786 22.441 59.548 22.515 ;
        RECT 52.74 22.487 59.502 22.561 ;
        RECT 52.694 22.533 59.456 22.607 ;
        RECT 52.648 22.579 59.41 22.653 ;
        RECT 52.602 22.625 59.364 22.699 ;
        RECT 52.556 22.671 59.318 22.745 ;
        RECT 52.51 22.717 59.272 22.791 ;
        RECT 52.464 22.763 59.226 22.837 ;
        RECT 52.418 22.809 59.18 22.883 ;
        RECT 52.372 22.855 59.134 22.929 ;
        RECT 52.326 22.901 59.088 22.975 ;
        RECT 52.28 22.947 59.042 23.021 ;
        RECT 52.234 22.993 58.996 23.067 ;
        RECT 52.188 23.039 58.95 23.113 ;
        RECT 52.142 23.085 58.904 23.159 ;
        RECT 52.096 23.131 58.858 23.205 ;
        RECT 52.05 23.177 58.812 23.251 ;
        RECT 52.004 23.223 58.766 23.297 ;
        RECT 51.958 23.269 58.72 23.343 ;
        RECT 51.912 23.315 58.674 23.389 ;
        RECT 51.866 23.361 58.628 23.435 ;
        RECT 51.82 23.407 58.582 23.481 ;
        RECT 51.774 23.453 58.536 23.527 ;
        RECT 51.728 23.499 58.49 23.573 ;
        RECT 51.682 23.545 58.444 23.619 ;
        RECT 51.636 23.591 58.398 23.665 ;
        RECT 51.59 23.637 58.352 23.711 ;
        RECT 51.544 23.683 58.306 23.757 ;
        RECT 51.498 23.729 58.26 23.803 ;
        RECT 51.452 23.775 58.214 23.849 ;
        RECT 51.406 23.821 58.168 23.895 ;
        RECT 51.36 23.867 58.122 23.941 ;
        RECT 51.314 23.913 58.076 23.987 ;
        RECT 51.268 23.959 58.03 24.033 ;
        RECT 51.222 24.005 57.984 24.079 ;
        RECT 51.176 24.051 57.938 24.125 ;
        RECT 51.13 24.097 57.892 24.171 ;
        RECT 51.084 24.143 57.846 24.217 ;
        RECT 51.038 24.189 57.8 24.263 ;
        RECT 50.992 24.235 57.754 24.309 ;
        RECT 50.946 24.281 57.708 24.355 ;
        RECT 50.9 24.327 57.662 24.401 ;
        RECT 50.854 24.373 57.616 24.447 ;
        RECT 50.808 24.419 57.57 24.493 ;
        RECT 50.762 24.465 57.524 24.539 ;
        RECT 50.716 24.511 57.478 24.585 ;
        RECT 50.67 24.557 57.432 24.631 ;
        RECT 50.624 24.603 57.386 24.677 ;
        RECT 50.578 24.649 57.34 24.723 ;
        RECT 50.532 24.695 57.294 24.769 ;
        RECT 50.486 24.741 57.248 24.815 ;
        RECT 50.44 24.787 57.202 24.861 ;
        RECT 50.394 24.833 57.156 24.907 ;
        RECT 50.348 24.879 57.11 24.953 ;
        RECT 50.302 24.925 57.064 24.999 ;
        RECT 50.256 24.971 57.018 25.045 ;
        RECT 50.21 25.017 56.972 25.091 ;
        RECT 50.164 25.063 56.926 25.137 ;
        RECT 50.118 25.109 56.88 25.183 ;
        RECT 50.072 25.155 56.834 25.229 ;
        RECT 50.026 25.201 56.788 25.275 ;
        RECT 49.98 25.247 56.742 25.321 ;
        RECT 49.934 25.293 56.696 25.367 ;
        RECT 49.888 25.339 56.65 25.413 ;
        RECT 49.842 25.385 56.604 25.459 ;
        RECT 49.796 25.431 56.558 25.505 ;
        RECT 49.75 25.477 56.512 25.551 ;
        RECT 49.704 25.523 56.466 25.597 ;
        RECT 49.658 25.569 56.42 25.643 ;
        RECT 49.612 25.615 56.374 25.689 ;
        RECT 49.566 25.661 56.328 25.735 ;
        RECT 49.52 25.707 56.282 25.781 ;
        RECT 49.474 25.753 56.236 25.827 ;
        RECT 49.428 25.799 56.19 25.873 ;
        RECT 49.382 25.845 56.144 25.919 ;
        RECT 49.336 25.891 56.098 25.965 ;
        RECT 49.29 25.937 56.052 26.011 ;
        RECT 49.244 25.983 56.006 26.057 ;
        RECT 49.198 26.029 55.96 26.103 ;
        RECT 49.152 26.075 55.914 26.149 ;
        RECT 49.106 26.121 55.868 26.195 ;
        RECT 49.06 26.167 55.822 26.241 ;
        RECT 49.014 26.213 55.776 26.287 ;
        RECT 48.968 26.259 55.73 26.333 ;
        RECT 48.922 26.305 55.684 26.379 ;
        RECT 48.876 26.351 55.638 26.425 ;
        RECT 48.83 26.397 55.592 26.471 ;
        RECT 48.784 26.443 55.546 26.517 ;
        RECT 48.738 26.489 55.5 26.563 ;
        RECT 48.692 26.535 55.454 26.609 ;
        RECT 48.646 26.581 55.408 26.655 ;
        RECT 48.6 26.627 55.362 26.701 ;
        RECT 48.554 26.673 55.316 26.747 ;
        RECT 48.508 26.719 55.27 26.793 ;
        RECT 48.462 26.765 55.224 26.839 ;
        RECT 48.416 26.811 55.178 26.885 ;
        RECT 48.37 26.857 55.132 26.931 ;
        RECT 48.324 26.903 55.086 26.977 ;
        RECT 48.278 26.949 55.04 27.023 ;
        RECT 48.232 26.995 54.994 27.069 ;
        RECT 48.186 27.041 54.948 27.115 ;
        RECT 48.14 27.087 54.902 27.161 ;
        RECT 48.094 27.133 54.856 27.207 ;
        RECT 48.048 27.179 54.81 27.253 ;
        RECT 48.002 27.225 54.764 27.299 ;
        RECT 47.956 27.271 54.718 27.345 ;
        RECT 47.91 27.317 54.672 27.391 ;
        RECT 47.864 27.363 54.626 27.437 ;
        RECT 47.818 27.409 54.58 27.483 ;
        RECT 47.772 27.455 54.534 27.529 ;
        RECT 47.726 27.501 54.488 27.575 ;
        RECT 47.68 27.547 54.442 27.621 ;
        RECT 47.634 27.593 54.396 27.667 ;
        RECT 47.588 27.639 54.35 27.713 ;
        RECT 47.542 27.685 54.304 27.759 ;
        RECT 47.496 27.731 54.258 27.805 ;
        RECT 47.45 27.777 54.212 27.851 ;
        RECT 47.404 27.823 54.166 27.897 ;
        RECT 47.358 27.869 54.12 27.943 ;
        RECT 47.312 27.915 54.074 27.989 ;
        RECT 47.266 27.961 54.028 28.035 ;
        RECT 47.22 28.007 53.982 28.081 ;
        RECT 47.174 28.053 53.936 28.127 ;
        RECT 47.128 28.099 53.89 28.173 ;
        RECT 47.082 28.145 53.844 28.219 ;
        RECT 47.036 28.191 53.798 28.265 ;
        RECT 46.99 28.237 53.752 28.311 ;
        RECT 46.944 28.283 53.706 28.357 ;
        RECT 46.898 28.329 53.66 28.403 ;
        RECT 46.852 28.375 53.614 28.449 ;
        RECT 46.806 28.421 53.568 28.495 ;
        RECT 46.76 28.467 53.522 28.541 ;
        RECT 46.714 28.513 53.476 28.587 ;
        RECT 46.668 28.559 53.43 28.633 ;
        RECT 46.622 28.605 53.384 28.679 ;
        RECT 46.576 28.651 53.338 28.725 ;
        RECT 46.53 28.697 53.292 28.771 ;
        RECT 46.484 28.743 53.246 28.817 ;
        RECT 46.438 28.789 53.2 28.863 ;
        RECT 46.392 28.835 53.154 28.909 ;
        RECT 46.346 28.881 53.108 28.955 ;
        RECT 46.3 28.927 53.062 29.001 ;
        RECT 46.254 28.973 53.016 29.047 ;
        RECT 46.208 29.019 52.97 29.093 ;
        RECT 46.162 29.065 52.924 29.139 ;
        RECT 46.116 29.111 52.878 29.185 ;
        RECT 46.07 29.157 52.832 29.231 ;
        RECT 46.024 29.203 52.786 29.277 ;
        RECT 45.978 29.249 52.74 29.323 ;
        RECT 45.932 29.295 52.694 29.369 ;
        RECT 45.886 29.341 52.648 29.415 ;
        RECT 45.84 29.387 52.602 29.461 ;
        RECT 45.794 29.433 52.556 29.507 ;
        RECT 45.748 29.479 52.51 29.553 ;
        RECT 45.702 29.525 52.464 29.599 ;
        RECT 45.656 29.571 52.418 29.645 ;
        RECT 45.61 29.617 52.372 29.691 ;
        RECT 45.564 29.663 52.326 29.737 ;
        RECT 45.518 29.709 52.28 29.783 ;
        RECT 45.472 29.755 52.234 29.829 ;
        RECT 45.426 29.801 52.188 29.875 ;
        RECT 45.38 29.847 52.142 29.921 ;
        RECT 45.334 29.893 52.096 29.967 ;
        RECT 45.288 29.939 52.05 30.013 ;
        RECT 45.242 29.985 52.004 30.059 ;
        RECT 45.196 30.031 51.958 30.105 ;
        RECT 45.15 30.077 51.912 30.151 ;
        RECT 45.104 30.123 51.866 30.197 ;
        RECT 45.058 30.169 51.82 30.243 ;
        RECT 45.012 30.215 51.774 30.289 ;
        RECT 44.966 30.261 51.728 30.335 ;
        RECT 44.92 30.307 51.682 30.381 ;
        RECT 44.874 30.353 51.636 30.427 ;
        RECT 44.828 30.399 51.59 30.473 ;
        RECT 44.782 30.445 51.544 30.519 ;
        RECT 44.736 30.491 51.498 30.565 ;
        RECT 44.69 30.537 51.452 30.611 ;
        RECT 44.644 30.583 51.406 30.657 ;
        RECT 44.598 30.629 51.36 30.703 ;
        RECT 44.552 30.675 51.314 30.749 ;
        RECT 44.506 30.721 51.268 30.795 ;
        RECT 44.46 30.767 51.222 30.841 ;
        RECT 44.414 30.813 51.176 30.887 ;
        RECT 44.368 30.859 51.13 30.933 ;
        RECT 44.322 30.905 51.084 30.979 ;
        RECT 44.276 30.951 51.038 31.025 ;
        RECT 44.23 30.997 50.992 31.071 ;
        RECT 44.184 31.043 50.946 31.117 ;
        RECT 44.138 31.089 50.9 31.163 ;
        RECT 44.092 31.135 50.854 31.209 ;
        RECT 44.046 31.181 50.808 31.255 ;
        RECT 44 31.227 50.762 31.301 ;
        RECT 43.954 31.273 50.716 31.347 ;
        RECT 43.908 31.319 50.67 31.393 ;
        RECT 43.862 31.365 50.624 31.439 ;
        RECT 43.816 31.411 50.578 31.485 ;
        RECT 43.77 31.457 50.532 31.531 ;
        RECT 43.724 31.503 50.486 31.577 ;
        RECT 43.678 31.549 50.44 31.623 ;
        RECT 43.632 31.595 50.394 31.669 ;
        RECT 43.586 31.641 50.348 31.715 ;
        RECT 43.54 31.687 50.302 31.761 ;
        RECT 43.494 31.733 50.256 31.807 ;
        RECT 43.448 31.779 50.21 31.853 ;
        RECT 43.402 31.825 50.164 31.899 ;
        RECT 43.356 31.871 50.118 31.945 ;
        RECT 43.31 31.917 50.072 31.991 ;
        RECT 43.264 31.963 50.026 32.037 ;
        RECT 43.218 32.009 49.98 32.083 ;
        RECT 43.172 32.055 49.934 32.129 ;
        RECT 43.126 32.101 49.888 32.175 ;
        RECT 43.08 32.147 49.842 32.221 ;
        RECT 43.034 32.193 49.796 32.267 ;
        RECT 42.988 32.239 49.75 32.313 ;
        RECT 42.942 32.285 49.704 32.359 ;
        RECT 42.896 32.331 49.658 32.405 ;
        RECT 42.85 32.377 49.612 32.451 ;
        RECT 42.804 32.423 49.566 32.497 ;
        RECT 42.758 32.469 49.52 32.543 ;
        RECT 42.712 32.515 49.474 32.589 ;
        RECT 42.666 32.561 49.428 32.635 ;
        RECT 42.62 32.607 49.382 32.681 ;
        RECT 42.574 32.653 49.336 32.727 ;
        RECT 42.528 32.699 49.29 32.773 ;
        RECT 42.482 32.745 49.244 32.819 ;
        RECT 42.436 32.791 49.198 32.865 ;
        RECT 42.39 32.837 49.152 32.911 ;
        RECT 42.344 32.883 49.106 32.957 ;
        RECT 42.298 32.929 49.06 33.003 ;
        RECT 42.252 32.975 49.014 33.049 ;
        RECT 42.206 33.021 48.968 33.095 ;
        RECT 42.16 33.067 48.922 33.141 ;
        RECT 42.114 33.113 48.876 33.187 ;
        RECT 42.068 33.159 48.83 33.233 ;
        RECT 42.022 33.205 48.784 33.279 ;
        RECT 41.976 33.251 48.738 33.325 ;
        RECT 41.93 33.297 48.692 33.371 ;
        RECT 41.884 33.343 48.646 33.417 ;
        RECT 41.838 33.389 48.6 33.463 ;
        RECT 41.792 33.435 48.554 33.509 ;
        RECT 41.746 33.481 48.508 33.555 ;
        RECT 41.7 33.527 48.462 33.601 ;
        RECT 41.654 33.573 48.416 33.647 ;
        RECT 41.608 33.619 48.37 33.693 ;
        RECT 41.562 33.665 48.324 33.739 ;
        RECT 41.516 33.711 48.278 33.785 ;
        RECT 41.47 33.757 48.232 33.831 ;
        RECT 41.424 33.803 48.186 33.877 ;
        RECT 41.378 33.849 48.14 33.923 ;
        RECT 41.332 33.895 48.094 33.969 ;
        RECT 41.286 33.941 48.048 34.015 ;
        RECT 41.24 33.987 48.002 34.061 ;
        RECT 41.194 34.033 47.956 34.107 ;
        RECT 41.148 34.079 47.91 34.153 ;
        RECT 41.102 34.125 47.864 34.199 ;
        RECT 41.056 34.171 47.818 34.245 ;
        RECT 41.01 34.217 47.772 34.291 ;
        RECT 40.964 34.263 47.726 34.337 ;
        RECT 40.918 34.309 47.68 34.383 ;
        RECT 40.872 34.355 47.634 34.429 ;
        RECT 40.826 34.401 47.588 34.475 ;
        RECT 40.78 34.447 47.542 34.521 ;
        RECT 40.734 34.493 47.496 34.567 ;
        RECT 40.688 34.539 47.45 34.613 ;
        RECT 40.642 34.585 47.404 34.659 ;
        RECT 40.596 34.631 47.358 34.705 ;
        RECT 40.55 34.677 47.312 34.751 ;
        RECT 40.504 34.723 47.266 34.797 ;
        RECT 40.458 34.769 47.22 34.843 ;
        RECT 40.412 34.815 47.174 34.889 ;
        RECT 40.366 34.861 47.128 34.935 ;
        RECT 40.32 34.907 47.082 34.981 ;
        RECT 40.274 34.953 47.036 35.027 ;
        RECT 40.228 34.999 46.99 35.073 ;
        RECT 40.182 35.045 46.944 35.119 ;
        RECT 40.136 35.091 46.898 35.165 ;
        RECT 40.09 35.137 46.852 35.211 ;
        RECT 40.044 35.183 46.806 35.257 ;
        RECT 39.998 35.229 46.76 35.303 ;
        RECT 39.952 35.275 46.714 35.349 ;
        RECT 39.906 35.321 46.668 35.395 ;
        RECT 39.86 35.367 46.622 35.441 ;
        RECT 39.814 35.413 46.576 35.487 ;
        RECT 39.768 35.459 46.53 35.533 ;
        RECT 39.722 35.505 46.484 35.579 ;
        RECT 39.676 35.551 46.438 35.625 ;
        RECT 39.63 35.597 46.392 35.671 ;
        RECT 39.584 35.643 46.346 35.717 ;
        RECT 39.538 35.689 46.3 35.763 ;
        RECT 39.492 35.735 46.254 35.809 ;
        RECT 39.446 35.781 46.208 35.855 ;
        RECT 39.4 35.827 46.162 35.901 ;
        RECT 39.354 35.873 46.116 35.947 ;
        RECT 39.308 35.919 46.07 35.993 ;
        RECT 39.262 35.965 46.024 36.039 ;
        RECT 39.216 36.011 45.978 36.085 ;
        RECT 39.17 36.057 45.932 36.131 ;
        RECT 39.124 36.103 45.886 36.177 ;
        RECT 39.078 36.149 45.84 36.223 ;
        RECT 39.032 36.195 45.794 36.269 ;
        RECT 38.986 36.241 45.748 36.315 ;
        RECT 38.94 36.287 45.702 36.361 ;
        RECT 38.894 36.333 45.656 36.407 ;
        RECT 38.848 36.379 45.61 36.453 ;
        RECT 38.802 36.425 45.564 36.499 ;
        RECT 38.756 36.471 45.518 36.545 ;
        RECT 38.71 36.517 45.472 36.591 ;
        RECT 38.664 36.563 45.426 36.637 ;
        RECT 38.618 36.609 45.38 36.683 ;
        RECT 38.572 36.655 45.334 36.729 ;
        RECT 38.526 36.701 45.288 36.775 ;
        RECT 38.48 36.747 45.242 36.821 ;
        RECT 38.434 36.793 45.196 36.867 ;
        RECT 38.388 36.839 45.15 36.913 ;
        RECT 38.342 36.885 45.104 36.959 ;
        RECT 38.296 36.931 45.058 37.005 ;
        RECT 38.25 36.977 45.012 37.051 ;
        RECT 38.204 37.023 44.966 37.097 ;
        RECT 38.158 37.069 44.92 37.143 ;
        RECT 38.112 37.115 44.874 37.189 ;
        RECT 38.066 37.161 44.828 37.235 ;
        RECT 38.02 37.207 44.782 37.281 ;
        RECT 37.974 37.253 44.736 37.327 ;
        RECT 37.928 37.299 44.69 37.373 ;
        RECT 37.882 37.345 44.644 37.419 ;
        RECT 37.836 37.391 44.598 37.465 ;
        RECT 37.79 37.437 44.552 37.511 ;
        RECT 37.744 37.483 44.506 37.557 ;
        RECT 37.698 37.529 44.46 37.603 ;
        RECT 37.652 37.575 44.414 37.649 ;
        RECT 37.606 37.621 44.368 37.695 ;
        RECT 37.56 37.667 44.322 37.741 ;
        RECT 37.514 37.713 44.276 37.787 ;
        RECT 37.468 37.759 44.23 37.833 ;
        RECT 37.422 37.805 44.184 37.879 ;
        RECT 37.376 37.851 44.138 37.925 ;
        RECT 37.33 37.897 44.092 37.971 ;
        RECT 37.284 37.943 44.046 38.017 ;
        RECT 37.238 37.989 44 38.063 ;
        RECT 37.192 38.035 43.954 38.109 ;
        RECT 37.146 38.081 43.908 38.155 ;
        RECT 37.1 38.127 43.862 38.201 ;
        RECT 37.054 38.173 43.816 38.247 ;
        RECT 37.008 38.219 43.77 38.293 ;
        RECT 36.962 38.265 43.724 38.339 ;
        RECT 36.916 38.311 43.678 38.385 ;
        RECT 36.87 38.357 43.632 38.431 ;
        RECT 36.824 38.403 43.586 38.477 ;
        RECT 36.778 38.449 43.54 38.523 ;
        RECT 36.732 38.495 43.494 38.569 ;
        RECT 36.686 38.541 43.448 38.615 ;
        RECT 36.64 38.587 43.402 38.661 ;
        RECT 36.594 38.633 43.356 38.707 ;
        RECT 36.548 38.679 43.31 38.753 ;
        RECT 36.502 38.725 43.264 38.799 ;
        RECT 36.456 38.771 43.218 38.845 ;
        RECT 36.41 38.817 43.172 38.891 ;
        RECT 36.364 38.863 43.126 38.937 ;
        RECT 36.318 38.909 43.08 38.983 ;
        RECT 36.272 38.955 43.034 39.029 ;
        RECT 36.226 39.001 42.988 39.075 ;
        RECT 36.18 39.047 42.942 39.121 ;
        RECT 36.134 39.093 42.896 39.167 ;
        RECT 36.088 39.139 42.85 39.213 ;
        RECT 36.042 39.185 42.804 39.259 ;
        RECT 35.996 39.231 42.758 39.305 ;
        RECT 35.95 39.277 42.712 39.351 ;
        RECT 35.904 39.323 42.666 39.397 ;
        RECT 35.858 39.369 42.62 39.443 ;
        RECT 35.812 39.415 42.574 39.489 ;
        RECT 35.766 39.461 42.528 39.535 ;
        RECT 35.72 39.507 42.482 39.581 ;
        RECT 35.674 39.553 42.436 39.627 ;
        RECT 35.628 39.599 42.39 39.673 ;
        RECT 35.582 39.645 42.344 39.719 ;
        RECT 35.536 39.691 42.298 39.765 ;
        RECT 35.49 39.737 42.252 39.811 ;
        RECT 35.444 39.783 42.206 39.857 ;
        RECT 35.398 39.829 42.16 39.903 ;
        RECT 35.352 39.875 42.114 39.949 ;
        RECT 35.306 39.921 42.068 39.995 ;
        RECT 35.26 39.967 42.022 40.041 ;
        RECT 35.214 40.013 41.976 40.087 ;
        RECT 35.168 40.059 41.93 40.133 ;
        RECT 35.122 40.105 41.884 40.179 ;
        RECT 35.076 40.151 41.838 40.225 ;
        RECT 35.03 40.197 41.792 40.271 ;
        RECT 34.984 40.243 41.746 40.317 ;
        RECT 34.938 40.289 41.7 40.363 ;
        RECT 34.892 40.335 41.654 40.409 ;
        RECT 34.846 40.381 41.608 40.455 ;
        RECT 34.8 40.427 41.562 40.501 ;
        RECT 34.754 40.473 41.516 40.547 ;
        RECT 34.708 40.519 41.47 40.593 ;
        RECT 34.662 40.565 41.424 40.639 ;
        RECT 34.616 40.611 41.378 40.685 ;
        RECT 34.57 40.657 41.332 40.731 ;
        RECT 34.524 40.703 41.286 40.777 ;
        RECT 34.478 40.749 41.24 40.823 ;
        RECT 34.432 40.795 41.194 40.869 ;
        RECT 34.386 40.841 41.148 40.915 ;
        RECT 34.34 40.887 41.102 40.961 ;
        RECT 34.294 40.933 41.056 41.007 ;
        RECT 34.248 40.979 41.01 41.053 ;
        RECT 34.202 41.025 40.964 41.099 ;
        RECT 34.156 41.071 40.918 41.145 ;
        RECT 34.11 41.117 40.872 41.191 ;
        RECT 34.064 41.163 40.826 41.237 ;
        RECT 34.018 41.209 40.78 41.283 ;
        RECT 33.972 41.255 40.734 41.329 ;
        RECT 33.926 41.301 40.688 41.375 ;
        RECT 33.88 41.347 40.642 41.421 ;
        RECT 33.834 41.393 40.596 41.467 ;
        RECT 33.788 41.439 40.55 41.513 ;
        RECT 33.742 41.485 40.504 41.559 ;
        RECT 33.696 41.531 40.458 41.605 ;
        RECT 33.65 41.577 40.412 41.651 ;
        RECT 33.604 41.623 40.366 41.697 ;
        RECT 33.558 41.669 40.32 41.743 ;
        RECT 33.512 41.715 40.274 41.789 ;
        RECT 33.466 41.761 40.228 41.835 ;
        RECT 33.42 41.807 40.182 41.881 ;
        RECT 33.374 41.853 40.136 41.927 ;
        RECT 33.328 41.899 40.09 41.973 ;
        RECT 33.282 41.945 40.044 42.019 ;
        RECT 33.236 41.991 39.998 42.065 ;
        RECT 33.19 42.037 39.952 42.111 ;
        RECT 33.144 42.083 39.906 42.157 ;
        RECT 33.098 42.129 39.86 42.203 ;
        RECT 33.052 42.175 39.814 42.249 ;
        RECT 33.006 42.221 39.768 42.295 ;
        RECT 32.96 42.267 39.722 42.341 ;
        RECT 32.914 42.313 39.676 42.387 ;
        RECT 32.868 42.359 39.63 42.433 ;
        RECT 32.822 42.405 39.584 42.479 ;
        RECT 32.776 42.451 39.538 42.525 ;
        RECT 32.73 42.497 39.492 42.571 ;
        RECT 32.684 42.543 39.446 42.617 ;
        RECT 32.638 42.589 39.4 42.663 ;
        RECT 32.592 42.635 39.354 42.709 ;
        RECT 32.546 42.681 39.308 42.755 ;
        RECT 32.5 42.727 39.262 42.801 ;
        RECT 32.454 42.773 39.216 42.847 ;
        RECT 32.408 42.819 39.17 42.893 ;
        RECT 32.362 42.865 39.124 42.939 ;
        RECT 32.316 42.911 39.078 42.985 ;
        RECT 32.27 42.957 39.032 43.031 ;
        RECT 32.224 43.003 38.986 43.077 ;
        RECT 32.178 43.049 38.94 43.123 ;
        RECT 32.132 43.095 38.894 43.169 ;
        RECT 32.086 43.141 38.848 43.215 ;
        RECT 32.04 43.187 38.802 43.261 ;
        RECT 31.994 43.233 38.756 43.307 ;
        RECT 31.948 43.279 38.71 43.353 ;
        RECT 31.902 43.325 38.664 43.399 ;
        RECT 31.856 43.371 38.618 43.445 ;
        RECT 31.81 43.417 38.572 43.491 ;
        RECT 31.764 43.463 38.526 43.537 ;
        RECT 31.718 43.509 38.48 43.583 ;
        RECT 31.672 43.555 38.434 43.629 ;
        RECT 31.626 43.601 38.388 43.675 ;
        RECT 31.58 43.647 38.342 43.721 ;
        RECT 31.534 43.693 38.296 43.767 ;
        RECT 31.488 43.739 38.25 43.813 ;
        RECT 31.442 43.785 38.204 43.859 ;
        RECT 31.396 43.831 38.158 43.905 ;
        RECT 31.35 43.877 38.112 43.951 ;
        RECT 31.304 43.923 38.066 43.997 ;
        RECT 31.258 43.969 38.02 44.043 ;
        RECT 31.212 44.015 37.974 44.089 ;
        RECT 31.166 44.061 37.928 44.135 ;
        RECT 31.12 44.107 37.882 44.181 ;
        RECT 31.074 44.153 37.836 44.227 ;
        RECT 31.028 44.199 37.79 44.273 ;
        RECT 30.982 44.245 37.744 44.319 ;
        RECT 30.936 44.291 37.698 44.365 ;
        RECT 30.89 44.337 37.652 44.411 ;
        RECT 30.844 44.383 37.606 44.457 ;
        RECT 30.798 44.429 37.56 44.503 ;
        RECT 30.752 44.475 37.514 44.549 ;
        RECT 30.706 44.521 37.468 44.595 ;
        RECT 30.66 44.567 37.422 44.641 ;
        RECT 30.614 44.613 37.376 44.687 ;
        RECT 30.568 44.659 37.33 44.733 ;
        RECT 30.522 44.705 37.284 44.779 ;
        RECT 30.476 44.751 37.238 44.825 ;
        RECT 30.43 44.797 37.192 44.871 ;
        RECT 30.384 44.843 37.146 44.917 ;
        RECT 30.338 44.889 37.1 44.963 ;
        RECT 30.292 44.935 37.054 45.009 ;
        RECT 30.246 44.981 37.008 45.055 ;
        RECT 30.2 45.027 36.962 45.101 ;
        RECT 30.154 45.073 36.916 45.147 ;
        RECT 30.108 45.119 36.87 45.193 ;
        RECT 30.062 45.165 36.824 45.239 ;
        RECT 30.016 45.211 36.778 45.285 ;
        RECT 29.97 45.257 36.732 45.331 ;
        RECT 29.924 45.303 36.686 45.377 ;
        RECT 29.878 45.349 36.64 45.423 ;
        RECT 29.832 45.395 36.594 45.469 ;
        RECT 29.786 45.441 36.548 45.515 ;
        RECT 29.74 45.487 36.502 45.561 ;
        RECT 29.694 45.533 36.456 45.607 ;
        RECT 29.648 45.579 36.41 45.653 ;
        RECT 29.602 45.625 36.364 45.699 ;
        RECT 29.556 45.671 36.318 45.745 ;
        RECT 29.51 45.717 36.272 45.791 ;
        RECT 29.464 45.763 36.226 45.837 ;
        RECT 29.418 45.809 36.18 45.883 ;
        RECT 29.372 45.855 36.134 45.929 ;
        RECT 29.326 45.901 36.088 45.975 ;
        RECT 29.28 45.947 36.042 46.021 ;
        RECT 29.234 45.993 35.996 46.067 ;
        RECT 29.188 46.039 35.95 46.113 ;
        RECT 29.142 46.085 35.904 46.159 ;
        RECT 29.096 46.131 35.858 46.205 ;
        RECT 29.05 46.177 35.812 46.251 ;
        RECT 29.004 46.223 35.766 46.297 ;
        RECT 28.958 46.269 35.72 46.343 ;
        RECT 28.912 46.315 35.674 46.389 ;
        RECT 28.866 46.361 35.628 46.435 ;
        RECT 28.82 46.407 35.582 46.481 ;
        RECT 28.774 46.453 35.536 46.527 ;
        RECT 28.728 46.499 35.49 46.573 ;
        RECT 28.682 46.545 35.444 46.619 ;
        RECT 28.636 46.591 35.398 46.665 ;
        RECT 28.59 46.637 35.352 46.711 ;
        RECT 28.544 46.683 35.306 46.757 ;
        RECT 28.498 46.729 35.26 46.803 ;
        RECT 28.452 46.775 35.214 46.849 ;
        RECT 28.406 46.821 35.168 46.895 ;
        RECT 28.36 46.867 35.122 46.941 ;
        RECT 28.314 46.913 35.076 46.987 ;
        RECT 28.268 46.959 35.03 47.033 ;
        RECT 28.222 47.005 34.984 47.079 ;
        RECT 28.176 47.051 34.938 47.125 ;
        RECT 28.13 47.097 34.892 47.171 ;
        RECT 28.084 47.143 34.846 47.217 ;
        RECT 28.038 47.189 34.8 47.263 ;
        RECT 27.992 47.235 34.754 47.309 ;
        RECT 27.946 47.281 34.708 47.355 ;
        RECT 27.9 47.327 34.662 47.401 ;
        RECT 27.854 47.373 34.616 47.447 ;
        RECT 27.808 47.419 34.57 47.493 ;
        RECT 27.762 47.465 34.524 47.539 ;
        RECT 27.716 47.511 34.478 47.585 ;
        RECT 27.67 47.557 34.432 47.631 ;
        RECT 27.624 47.603 34.386 47.677 ;
        RECT 27.578 47.649 34.34 47.723 ;
        RECT 27.532 47.695 34.294 47.769 ;
        RECT 27.486 47.741 34.248 47.815 ;
        RECT 27.44 47.787 34.202 47.861 ;
        RECT 27.394 47.833 34.156 47.907 ;
        RECT 27.348 47.879 34.11 47.953 ;
        RECT 27.302 47.925 34.064 47.999 ;
        RECT 27.256 47.971 34.018 48.045 ;
        RECT 27.21 48.017 33.972 48.091 ;
        RECT 27.164 48.063 33.926 48.137 ;
        RECT 27.118 48.109 33.88 48.183 ;
        RECT 27.072 48.155 33.834 48.229 ;
        RECT 27.026 48.201 33.788 48.275 ;
        RECT 26.98 48.247 33.742 48.321 ;
        RECT 26.934 48.293 33.696 48.367 ;
        RECT 26.888 48.339 33.65 48.413 ;
        RECT 26.842 48.385 33.604 48.459 ;
        RECT 26.796 48.431 33.558 48.505 ;
        RECT 26.75 48.477 33.512 48.551 ;
        RECT 26.704 48.523 33.466 48.597 ;
        RECT 26.658 48.569 33.42 48.643 ;
        RECT 26.612 48.615 33.374 48.689 ;
        RECT 26.566 48.661 33.328 48.735 ;
        RECT 26.52 48.707 33.282 48.781 ;
        RECT 26.474 48.753 33.236 48.827 ;
        RECT 26.428 48.799 33.19 48.873 ;
        RECT 26.382 48.845 33.144 48.919 ;
        RECT 26.336 48.891 33.098 48.965 ;
        RECT 26.29 48.937 33.052 49.011 ;
        RECT 26.244 48.983 33.006 49.057 ;
        RECT 26.198 49.029 32.96 49.103 ;
        RECT 26.152 49.075 32.914 49.149 ;
        RECT 26.106 49.121 32.868 49.195 ;
        RECT 26.06 49.167 32.822 49.241 ;
        RECT 26.014 49.213 32.776 49.287 ;
        RECT 25.968 49.259 32.73 49.333 ;
        RECT 25.922 49.305 32.684 49.379 ;
        RECT 25.876 49.351 32.638 49.425 ;
        RECT 25.83 49.397 32.592 49.471 ;
        RECT 25.784 49.443 32.546 49.517 ;
        RECT 25.738 49.489 32.5 49.563 ;
        RECT 25.692 49.535 32.454 49.609 ;
        RECT 25.646 49.581 32.408 49.655 ;
        RECT 25.6 49.627 32.362 49.701 ;
        RECT 25.554 49.673 32.316 49.747 ;
        RECT 25.508 49.719 32.27 49.793 ;
        RECT 25.462 49.765 32.224 49.839 ;
        RECT 25.416 49.811 32.178 49.885 ;
        RECT 25.37 49.857 32.132 49.931 ;
        RECT 25.324 49.903 32.086 49.977 ;
        RECT 25.278 49.949 32.04 50.023 ;
        RECT 25.232 49.995 31.994 50.069 ;
        RECT 25.186 50.041 31.948 50.115 ;
        RECT 25.14 50.087 31.902 50.161 ;
        RECT 25.094 50.133 31.856 50.207 ;
        RECT 25.048 50.179 31.81 50.253 ;
        RECT 25.002 50.225 31.764 50.299 ;
        RECT 24.956 50.271 31.718 50.345 ;
        RECT 24.91 50.317 31.672 50.391 ;
        RECT 24.864 50.363 31.626 50.437 ;
        RECT 24.818 50.409 31.58 50.483 ;
        RECT 24.772 50.455 31.534 50.529 ;
        RECT 24.726 50.501 31.488 50.575 ;
        RECT 24.68 50.547 31.442 50.621 ;
        RECT 24.634 50.593 31.396 50.667 ;
        RECT 24.588 50.639 31.35 50.713 ;
        RECT 24.542 50.685 31.304 50.759 ;
        RECT 24.496 50.731 31.258 50.805 ;
        RECT 24.45 50.777 31.212 50.851 ;
        RECT 24.404 50.823 31.166 50.897 ;
        RECT 24.358 50.869 31.12 50.943 ;
        RECT 24.312 50.915 31.074 50.989 ;
        RECT 24.266 50.961 31.028 51.035 ;
        RECT 24.22 51.007 30.982 51.081 ;
        RECT 24.174 51.053 30.936 51.127 ;
        RECT 24.128 51.099 30.89 51.173 ;
        RECT 24.082 51.145 30.844 51.219 ;
        RECT 24.036 51.191 30.798 51.265 ;
        RECT 23.99 51.237 30.752 51.311 ;
        RECT 23.944 51.283 30.706 51.357 ;
        RECT 23.898 51.329 30.66 51.403 ;
        RECT 23.852 51.375 30.614 51.449 ;
        RECT 23.806 51.421 30.568 51.495 ;
        RECT 23.76 51.467 30.522 51.541 ;
        RECT 23.714 51.513 30.476 51.587 ;
        RECT 23.668 51.559 30.43 51.633 ;
        RECT 23.622 51.605 30.384 51.679 ;
        RECT 23.576 51.651 30.338 51.725 ;
        RECT 23.53 51.697 30.292 51.771 ;
        RECT 23.484 51.743 30.246 51.817 ;
        RECT 23.438 51.789 30.2 51.863 ;
        RECT 23.392 51.835 30.154 51.909 ;
        RECT 23.346 51.881 30.108 51.955 ;
        RECT 23.3 51.927 30.062 52.001 ;
        RECT 23.254 51.973 30.016 52.047 ;
        RECT 23.208 52.019 29.97 52.093 ;
        RECT 23.162 52.065 29.924 52.139 ;
        RECT 23.116 52.111 29.878 52.185 ;
        RECT 23.07 52.157 29.832 52.231 ;
        RECT 23.024 52.203 29.786 52.277 ;
        RECT 22.978 52.249 29.74 52.323 ;
        RECT 22.932 52.295 29.694 52.369 ;
        RECT 22.886 52.341 29.648 52.415 ;
        RECT 22.84 52.387 29.602 52.461 ;
        RECT 22.794 52.433 29.556 52.507 ;
        RECT 22.748 52.479 29.51 52.553 ;
        RECT 22.702 52.525 29.464 52.599 ;
        RECT 22.656 52.571 29.418 52.645 ;
        RECT 22.61 52.617 29.372 52.691 ;
        RECT 22.564 52.663 29.326 52.737 ;
        RECT 22.518 52.709 29.28 52.783 ;
        RECT 22.472 52.755 29.234 52.829 ;
        RECT 22.426 52.801 29.188 52.875 ;
        RECT 22.38 52.847 29.142 52.921 ;
        RECT 22.334 52.893 29.096 52.967 ;
        RECT 22.288 52.939 29.05 53.013 ;
        RECT 22.242 52.985 29.004 53.059 ;
        RECT 22.196 53.031 28.958 53.105 ;
        RECT 22.15 53.077 28.912 53.151 ;
        RECT 22.104 53.123 28.866 53.197 ;
        RECT 22.058 53.169 28.82 53.243 ;
        RECT 22.012 53.215 28.774 53.289 ;
        RECT 21.966 53.261 28.728 53.335 ;
        RECT 21.92 53.307 28.682 53.381 ;
        RECT 21.874 53.353 28.636 53.427 ;
        RECT 21.828 53.399 28.59 53.473 ;
        RECT 21.782 53.445 28.544 53.519 ;
        RECT 21.736 53.491 28.498 53.565 ;
        RECT 21.69 53.537 28.452 53.611 ;
        RECT 21.644 53.583 28.406 53.657 ;
        RECT 21.598 53.629 28.36 53.703 ;
        RECT 21.552 53.675 28.314 53.749 ;
        RECT 21.506 53.721 28.268 53.795 ;
        RECT 21.46 53.767 28.222 53.841 ;
        RECT 21.414 53.813 28.176 53.887 ;
        RECT 21.368 53.859 28.13 53.933 ;
        RECT 21.322 53.905 28.084 53.979 ;
        RECT 21.276 53.951 28.038 54.025 ;
        RECT 21.23 53.997 27.992 54.071 ;
        RECT 21.184 54.043 27.946 54.117 ;
        RECT 21.138 54.089 27.9 54.163 ;
        RECT 21.092 54.135 27.854 54.209 ;
        RECT 21.046 54.181 27.808 54.255 ;
        RECT 21 54.227 27.762 54.301 ;
        RECT 20.954 54.273 27.716 54.347 ;
        RECT 20.908 54.319 27.67 54.393 ;
        RECT 20.862 54.365 27.624 54.439 ;
        RECT 20.816 54.411 27.578 54.485 ;
        RECT 20.77 54.457 27.532 54.531 ;
        RECT 20.724 54.503 27.486 54.577 ;
        RECT 20.678 54.549 27.44 54.623 ;
        RECT 20.632 54.595 27.394 54.669 ;
        RECT 20.586 54.641 27.348 54.715 ;
        RECT 20.54 54.687 27.302 54.761 ;
        RECT 20.494 54.733 27.256 54.807 ;
        RECT 20.448 54.779 27.21 54.853 ;
        RECT 20.402 54.825 27.164 54.899 ;
        RECT 20.356 54.871 27.118 54.945 ;
        RECT 20.31 54.917 27.072 54.991 ;
        RECT 20.264 54.963 27.026 55.037 ;
        RECT 20.218 55.009 26.98 55.083 ;
        RECT 20.172 55.055 26.934 55.129 ;
        RECT 20.126 55.101 26.888 55.175 ;
        RECT 20.08 55.147 26.842 55.221 ;
        RECT 20.034 55.193 26.796 55.267 ;
        RECT 19.988 55.239 26.75 55.313 ;
        RECT 19.942 55.285 26.704 55.359 ;
        RECT 19.896 55.331 26.658 55.405 ;
        RECT 19.85 55.377 26.612 55.451 ;
        RECT 19.804 55.423 26.566 55.497 ;
        RECT 19.758 55.469 26.52 55.543 ;
        RECT 19.712 55.515 26.474 55.589 ;
        RECT 19.666 55.561 26.428 55.635 ;
        RECT 19.62 55.607 26.382 55.681 ;
        RECT 19.574 55.653 26.336 55.727 ;
        RECT 19.528 55.699 26.29 55.773 ;
        RECT 19.482 55.745 26.244 55.819 ;
        RECT 19.436 55.791 26.198 55.865 ;
        RECT 19.39 55.837 26.152 55.911 ;
        RECT 19.344 55.883 26.106 55.957 ;
        RECT 19.298 55.929 26.06 56.003 ;
        RECT 19.252 55.975 26.014 56.049 ;
        RECT 19.206 56.021 25.968 56.095 ;
        RECT 19.16 56.067 25.922 56.141 ;
        RECT 19.114 56.113 25.876 56.187 ;
        RECT 19.068 56.159 25.83 56.233 ;
        RECT 19.022 56.205 25.784 56.279 ;
        RECT 18.976 56.251 25.738 56.325 ;
        RECT 18.93 56.297 25.692 56.371 ;
        RECT 18.884 56.343 25.646 56.417 ;
        RECT 18.838 56.389 25.6 56.463 ;
        RECT 18.792 56.435 25.554 56.509 ;
        RECT 18.746 56.481 25.508 56.555 ;
        RECT 18.7 56.527 25.462 56.601 ;
        RECT 18.654 56.573 25.416 56.647 ;
        RECT 18.608 56.619 25.37 56.693 ;
        RECT 18.562 56.665 25.324 56.739 ;
        RECT 18.516 56.711 25.278 56.785 ;
        RECT 18.47 56.757 25.232 56.831 ;
        RECT 18.424 56.803 25.186 56.877 ;
        RECT 18.378 56.849 25.14 56.923 ;
        RECT 18.332 56.895 25.094 56.969 ;
        RECT 18.286 56.941 25.048 57.015 ;
        RECT 18.24 56.987 25.002 57.061 ;
        RECT 18.194 57.033 24.956 57.107 ;
        RECT 18.148 57.079 24.91 57.153 ;
        RECT 18.102 57.125 24.864 57.199 ;
        RECT 18.056 57.171 24.818 57.245 ;
        RECT 18.01 57.217 24.772 57.291 ;
        RECT 17.964 57.263 24.726 57.337 ;
        RECT 17.918 57.309 24.68 57.383 ;
        RECT 17.872 57.355 24.634 57.429 ;
        RECT 17.826 57.401 24.588 57.475 ;
        RECT 17.78 57.447 24.542 57.521 ;
    END
    PORT
      LAYER QB ;
        RECT 59.462 42.075 66.218 42.155 ;
        RECT 64.108 37.429 64.154 44.219 ;
        RECT 57.346 44.191 64.108 44.265 ;
        RECT 59.508 42.029 66.264 42.109 ;
        RECT 64.062 37.475 64.108 44.265 ;
        RECT 57.3 44.237 64.062 44.311 ;
        RECT 59.554 41.983 66.31 42.063 ;
        RECT 64.016 37.521 64.062 44.311 ;
        RECT 57.254 44.283 64.016 44.357 ;
        RECT 59.6 41.937 66.356 42.017 ;
        RECT 63.97 37.567 64.016 44.357 ;
        RECT 57.208 44.329 63.97 44.403 ;
        RECT 59.646 41.891 66.402 41.971 ;
        RECT 63.924 37.613 63.97 44.403 ;
        RECT 57.162 44.375 63.924 44.449 ;
        RECT 59.692 41.845 66.448 41.925 ;
        RECT 63.878 37.659 63.924 44.449 ;
        RECT 57.116 44.421 63.878 44.495 ;
        RECT 59.738 41.799 66.494 41.879 ;
        RECT 63.832 37.705 63.878 44.495 ;
        RECT 57.07 44.467 63.832 44.541 ;
        RECT 59.784 41.753 66.54 41.833 ;
        RECT 63.786 37.751 63.832 44.541 ;
        RECT 57.024 44.513 63.786 44.587 ;
        RECT 59.83 41.707 66.586 41.787 ;
        RECT 63.74 37.797 63.786 44.587 ;
        RECT 56.978 44.559 63.74 44.633 ;
        RECT 59.876 41.661 66.632 41.741 ;
        RECT 63.694 37.843 63.74 44.633 ;
        RECT 56.932 44.605 63.694 44.679 ;
        RECT 59.922 41.615 66.678 41.695 ;
        RECT 63.648 37.889 63.694 44.679 ;
        RECT 56.886 44.651 63.648 44.725 ;
        RECT 59.968 41.569 66.724 41.649 ;
        RECT 63.602 37.935 63.648 44.725 ;
        RECT 56.84 44.697 63.602 44.771 ;
        RECT 60.014 41.523 66.77 41.603 ;
        RECT 63.556 37.981 63.602 44.771 ;
        RECT 56.794 44.743 63.556 44.817 ;
        RECT 60.06 41.477 66.816 41.557 ;
        RECT 63.51 38.027 63.556 44.817 ;
        RECT 56.748 44.789 63.51 44.863 ;
        RECT 60.106 41.431 66.862 41.511 ;
        RECT 63.464 38.073 63.51 44.863 ;
        RECT 56.702 44.835 63.464 44.909 ;
        RECT 60.152 41.385 66.908 41.465 ;
        RECT 63.418 38.119 63.464 44.909 ;
        RECT 56.656 44.881 63.418 44.955 ;
        RECT 60.198 41.339 66.954 41.419 ;
        RECT 63.372 38.165 63.418 44.955 ;
        RECT 56.61 44.927 63.372 45.001 ;
        RECT 60.244 41.293 67 41.373 ;
        RECT 63.326 38.211 63.372 45.001 ;
        RECT 56.564 44.973 63.326 45.047 ;
        RECT 60.29 41.247 67.046 41.327 ;
        RECT 63.28 38.257 63.326 45.047 ;
        RECT 56.518 45.019 63.28 45.093 ;
        RECT 60.336 41.201 67.092 41.281 ;
        RECT 63.234 38.303 63.28 45.093 ;
        RECT 56.472 45.065 63.234 45.139 ;
        RECT 60.428 41.109 80 41.2 ;
        RECT 63.188 38.349 63.234 45.139 ;
        RECT 56.426 45.111 63.188 45.185 ;
        RECT 60.474 41.063 80 41.2 ;
        RECT 63.142 38.395 63.188 45.185 ;
        RECT 56.38 45.157 63.142 45.231 ;
        RECT 60.52 41.017 80 41.2 ;
        RECT 63.096 38.441 63.142 45.231 ;
        RECT 56.334 45.203 63.096 45.277 ;
        RECT 60.566 40.971 80 41.2 ;
        RECT 63.05 38.487 63.096 45.277 ;
        RECT 56.288 45.249 63.05 45.323 ;
        RECT 60.612 40.925 80 41.2 ;
        RECT 63.004 38.533 63.05 45.323 ;
        RECT 56.242 45.295 63.004 45.369 ;
        RECT 60.658 40.879 80 41.2 ;
        RECT 62.958 38.579 63.004 45.369 ;
        RECT 56.196 45.341 62.958 45.415 ;
        RECT 60.704 40.833 80 41.2 ;
        RECT 62.912 38.625 62.958 45.415 ;
        RECT 56.15 45.387 62.912 45.461 ;
        RECT 60.75 40.787 80 41.2 ;
        RECT 62.866 38.671 62.912 45.461 ;
        RECT 56.104 45.433 62.866 45.507 ;
        RECT 60.796 40.741 80 41.2 ;
        RECT 62.82 38.717 62.866 45.507 ;
        RECT 56.058 45.479 62.82 45.553 ;
        RECT 60.842 40.695 80 41.2 ;
        RECT 62.774 38.763 62.82 45.553 ;
        RECT 56.012 45.525 62.774 45.599 ;
        RECT 60.888 40.649 80 41.2 ;
        RECT 62.728 38.809 62.774 45.599 ;
        RECT 55.966 45.571 62.728 45.645 ;
        RECT 60.934 40.603 80 41.2 ;
        RECT 62.682 38.855 62.728 45.645 ;
        RECT 55.92 45.617 62.682 45.691 ;
        RECT 60.98 40.557 80 41.2 ;
        RECT 62.636 38.901 62.682 45.691 ;
        RECT 55.874 45.663 62.636 45.737 ;
        RECT 61.026 40.511 80 41.2 ;
        RECT 62.59 38.947 62.636 45.737 ;
        RECT 55.828 45.709 62.59 45.783 ;
        RECT 61.072 40.465 80 41.2 ;
        RECT 62.544 38.993 62.59 45.783 ;
        RECT 55.782 45.755 62.544 45.829 ;
        RECT 61.118 40.419 80 41.2 ;
        RECT 62.498 39.039 62.544 45.829 ;
        RECT 55.736 45.801 62.498 45.875 ;
        RECT 61.164 40.373 80 41.2 ;
        RECT 62.452 39.085 62.498 45.875 ;
        RECT 55.69 45.847 62.452 45.921 ;
        RECT 61.21 40.327 80 41.2 ;
        RECT 62.406 39.131 62.452 45.921 ;
        RECT 55.644 45.893 62.406 45.967 ;
        RECT 61.256 40.281 80 41.2 ;
        RECT 62.36 39.177 62.406 45.967 ;
        RECT 55.598 45.939 62.36 46.013 ;
        RECT 61.302 40.235 80 41.2 ;
        RECT 62.314 39.223 62.36 46.013 ;
        RECT 55.552 45.985 62.314 46.059 ;
        RECT 61.348 40.189 80 41.2 ;
        RECT 62.268 39.269 62.314 46.059 ;
        RECT 55.506 46.031 62.268 46.105 ;
        RECT 61.394 40.143 80 41.2 ;
        RECT 62.222 39.315 62.268 46.105 ;
        RECT 55.46 46.077 62.222 46.151 ;
        RECT 61.44 40.097 80 41.2 ;
        RECT 62.176 39.361 62.222 46.151 ;
        RECT 55.414 46.123 62.176 46.197 ;
        RECT 61.486 40.051 80 41.2 ;
        RECT 62.13 39.407 62.176 46.197 ;
        RECT 55.368 46.169 62.13 46.243 ;
        RECT 61.532 40.005 80 41.2 ;
        RECT 62.084 39.453 62.13 46.243 ;
        RECT 55.322 46.215 62.084 46.289 ;
        RECT 61.578 39.959 80 41.2 ;
        RECT 62.038 39.499 62.084 46.289 ;
        RECT 55.276 46.261 62.038 46.335 ;
        RECT 61.624 39.913 80 41.2 ;
        RECT 61.992 39.545 62.038 46.335 ;
        RECT 55.23 46.307 61.992 46.381 ;
        RECT 61.67 39.867 80 41.2 ;
        RECT 61.946 39.591 61.992 46.381 ;
        RECT 55.184 46.353 61.946 46.427 ;
        RECT 61.716 39.821 80 41.2 ;
        RECT 61.9 39.637 61.946 46.427 ;
        RECT 55.138 46.399 61.9 46.473 ;
        RECT 61.762 39.775 80 41.2 ;
        RECT 61.854 39.683 61.9 46.473 ;
        RECT 55.092 46.445 61.854 46.519 ;
        RECT 61.808 39.729 80 41.2 ;
        RECT 55.046 46.491 61.808 46.565 ;
        RECT 55 46.537 61.762 46.611 ;
        RECT 54.954 46.583 61.716 46.657 ;
        RECT 54.908 46.629 61.67 46.703 ;
        RECT 54.862 46.675 61.624 46.749 ;
        RECT 54.816 46.721 61.578 46.795 ;
        RECT 54.77 46.767 61.532 46.841 ;
        RECT 54.724 46.813 61.486 46.887 ;
        RECT 54.678 46.859 61.44 46.933 ;
        RECT 54.632 46.905 61.394 46.979 ;
        RECT 54.586 46.951 61.348 47.025 ;
        RECT 54.54 46.997 61.302 47.071 ;
        RECT 54.494 47.043 61.256 47.117 ;
        RECT 54.448 47.089 61.21 47.163 ;
        RECT 54.402 47.135 61.164 47.209 ;
        RECT 54.356 47.181 61.118 47.255 ;
        RECT 54.31 47.227 61.072 47.301 ;
        RECT 54.264 47.273 61.026 47.347 ;
        RECT 54.218 47.319 60.98 47.393 ;
        RECT 54.172 47.365 60.934 47.439 ;
        RECT 54.126 47.411 60.888 47.485 ;
        RECT 54.08 47.457 60.842 47.531 ;
        RECT 54.034 47.503 60.796 47.577 ;
        RECT 53.988 47.549 60.75 47.623 ;
        RECT 53.942 47.595 60.704 47.669 ;
        RECT 53.896 47.641 60.658 47.715 ;
        RECT 53.85 47.687 60.612 47.761 ;
        RECT 53.804 47.733 60.566 47.807 ;
        RECT 53.758 47.779 60.52 47.853 ;
        RECT 53.712 47.825 60.474 47.899 ;
        RECT 53.666 47.871 60.428 47.945 ;
        RECT 53.62 47.917 60.382 47.991 ;
        RECT 53.574 47.963 60.336 48.037 ;
        RECT 53.528 48.009 60.29 48.083 ;
        RECT 53.482 48.055 60.244 48.129 ;
        RECT 53.436 48.101 60.198 48.175 ;
        RECT 53.39 48.147 60.152 48.221 ;
        RECT 53.344 48.193 60.106 48.267 ;
        RECT 53.298 48.239 60.06 48.313 ;
        RECT 53.252 48.285 60.014 48.359 ;
        RECT 53.206 48.331 59.968 48.405 ;
        RECT 53.16 48.377 59.922 48.451 ;
        RECT 53.114 48.423 59.876 48.497 ;
        RECT 53.068 48.469 59.83 48.543 ;
        RECT 53.022 48.515 59.784 48.589 ;
        RECT 52.976 48.561 59.738 48.635 ;
        RECT 52.93 48.607 59.692 48.681 ;
        RECT 52.884 48.653 59.646 48.727 ;
        RECT 52.838 48.699 59.6 48.773 ;
        RECT 52.792 48.745 59.554 48.819 ;
        RECT 52.746 48.791 59.508 48.865 ;
        RECT 52.7 48.837 59.462 48.911 ;
        RECT 52.654 48.883 59.416 48.957 ;
        RECT 52.608 48.929 59.37 49.003 ;
        RECT 52.562 48.975 59.324 49.049 ;
        RECT 52.516 49.021 59.278 49.095 ;
        RECT 52.47 49.067 59.232 49.141 ;
        RECT 52.424 49.113 59.186 49.187 ;
        RECT 52.378 49.159 59.14 49.233 ;
        RECT 52.332 49.205 59.094 49.279 ;
        RECT 52.286 49.251 59.048 49.325 ;
        RECT 52.24 49.297 59.002 49.371 ;
        RECT 52.194 49.343 58.956 49.417 ;
        RECT 52.148 49.389 58.91 49.463 ;
        RECT 52.102 49.435 58.864 49.509 ;
        RECT 52.056 49.481 58.818 49.555 ;
        RECT 52.01 49.527 58.772 49.601 ;
        RECT 51.964 49.573 58.726 49.647 ;
        RECT 51.918 49.619 58.68 49.693 ;
        RECT 51.872 49.665 58.634 49.739 ;
        RECT 51.826 49.711 58.588 49.785 ;
        RECT 51.78 49.757 58.542 49.831 ;
        RECT 51.734 49.803 58.496 49.877 ;
        RECT 51.688 49.849 58.45 49.923 ;
        RECT 51.642 49.895 58.404 49.969 ;
        RECT 51.596 49.941 58.358 50.015 ;
        RECT 51.55 49.987 58.312 50.061 ;
        RECT 51.504 50.033 58.266 50.107 ;
        RECT 51.458 50.079 58.22 50.153 ;
        RECT 51.412 50.125 58.174 50.199 ;
        RECT 51.366 50.171 58.128 50.245 ;
        RECT 51.32 50.217 58.082 50.291 ;
        RECT 51.274 50.263 58.036 50.337 ;
        RECT 51.228 50.309 57.99 50.383 ;
        RECT 51.182 50.355 57.944 50.429 ;
        RECT 51.136 50.401 57.898 50.475 ;
        RECT 51.09 50.447 57.852 50.521 ;
        RECT 51.044 50.493 57.806 50.567 ;
        RECT 50.998 50.539 57.76 50.613 ;
        RECT 50.952 50.585 57.714 50.659 ;
        RECT 50.906 50.631 57.668 50.705 ;
        RECT 50.86 50.677 57.622 50.751 ;
        RECT 50.814 50.723 57.576 50.797 ;
        RECT 50.768 50.769 57.53 50.843 ;
        RECT 50.722 50.815 57.484 50.889 ;
        RECT 50.676 50.861 57.438 50.935 ;
        RECT 50.63 50.907 57.392 50.981 ;
        RECT 50.584 50.953 57.346 51.027 ;
        RECT 50.538 50.999 57.3 51.073 ;
        RECT 50.492 51.045 57.254 51.119 ;
        RECT 50.446 51.091 57.208 51.165 ;
        RECT 50.4 51.137 57.162 51.211 ;
        RECT 50.354 51.183 57.116 51.257 ;
        RECT 50.308 51.229 57.07 51.303 ;
        RECT 50.262 51.275 57.024 51.349 ;
        RECT 50.216 51.321 56.978 51.395 ;
        RECT 50.17 51.367 56.932 51.441 ;
        RECT 50.124 51.413 56.886 51.487 ;
        RECT 50.078 51.459 56.84 51.533 ;
        RECT 50.032 51.505 56.794 51.579 ;
        RECT 49.986 51.551 56.748 51.625 ;
        RECT 49.94 51.597 56.702 51.671 ;
        RECT 49.894 51.643 56.656 51.717 ;
        RECT 49.848 51.689 56.61 51.763 ;
        RECT 49.802 51.735 56.564 51.809 ;
        RECT 49.756 51.781 56.518 51.855 ;
        RECT 49.71 51.827 56.472 51.901 ;
        RECT 49.664 51.873 56.426 51.947 ;
        RECT 49.618 51.919 56.38 51.993 ;
        RECT 49.572 51.965 56.334 52.039 ;
        RECT 49.526 52.011 56.288 52.085 ;
        RECT 49.48 52.057 56.242 52.131 ;
        RECT 49.434 52.103 56.196 52.177 ;
        RECT 49.388 52.149 56.15 52.223 ;
        RECT 49.342 52.195 56.104 52.269 ;
        RECT 49.296 52.241 56.058 52.315 ;
        RECT 49.25 52.287 56.012 52.361 ;
        RECT 49.204 52.333 55.966 52.407 ;
        RECT 49.158 52.379 55.92 52.453 ;
        RECT 49.112 52.425 55.874 52.499 ;
        RECT 49.066 52.471 55.828 52.545 ;
        RECT 49.02 52.517 55.782 52.591 ;
        RECT 48.974 52.563 55.736 52.637 ;
        RECT 48.928 52.609 55.69 52.683 ;
        RECT 48.882 52.655 55.644 52.729 ;
        RECT 48.836 52.701 55.598 52.775 ;
        RECT 48.79 52.747 55.552 52.821 ;
        RECT 48.744 52.793 55.506 52.867 ;
        RECT 48.698 52.839 55.46 52.913 ;
        RECT 48.652 52.885 55.414 52.959 ;
        RECT 48.606 52.931 55.368 53.005 ;
        RECT 48.56 52.977 55.322 53.051 ;
        RECT 48.514 53.023 55.276 53.097 ;
        RECT 48.468 53.069 55.23 53.143 ;
        RECT 48.422 53.115 55.184 53.189 ;
        RECT 48.376 53.161 55.138 53.235 ;
        RECT 48.33 53.207 55.092 53.281 ;
        RECT 48.284 53.253 55.046 53.327 ;
        RECT 48.238 53.299 55 53.373 ;
        RECT 48.192 53.345 54.954 53.419 ;
        RECT 48.146 53.391 54.908 53.465 ;
        RECT 48.1 53.437 54.862 53.511 ;
        RECT 48.054 53.483 54.816 53.557 ;
        RECT 48.008 53.529 54.77 53.603 ;
        RECT 47.962 53.575 54.724 53.649 ;
        RECT 47.916 53.621 54.678 53.695 ;
        RECT 47.87 53.667 54.632 53.741 ;
        RECT 47.824 53.713 54.586 53.787 ;
        RECT 47.778 53.759 54.54 53.833 ;
        RECT 47.732 53.805 54.494 53.879 ;
        RECT 47.686 53.851 54.448 53.925 ;
        RECT 47.64 53.897 54.402 53.971 ;
        RECT 47.594 53.943 54.356 54.017 ;
        RECT 47.548 53.989 54.31 54.063 ;
        RECT 47.502 54.035 54.264 54.109 ;
        RECT 47.456 54.081 54.218 54.155 ;
        RECT 47.41 54.127 54.172 54.201 ;
        RECT 47.364 54.173 54.126 54.247 ;
        RECT 47.318 54.219 54.08 54.293 ;
        RECT 47.272 54.265 54.034 54.339 ;
        RECT 47.226 54.311 53.988 54.385 ;
        RECT 47.18 54.357 53.942 54.431 ;
        RECT 47.134 54.403 53.896 54.477 ;
        RECT 47.088 54.449 53.85 54.523 ;
        RECT 47.042 54.495 53.804 54.569 ;
        RECT 46.996 54.541 53.758 54.615 ;
        RECT 46.95 54.587 53.712 54.661 ;
        RECT 46.904 54.633 53.666 54.707 ;
        RECT 46.858 54.679 53.62 54.753 ;
        RECT 46.812 54.725 53.574 54.799 ;
        RECT 46.766 54.771 53.528 54.845 ;
        RECT 46.72 54.817 53.482 54.891 ;
        RECT 46.674 54.863 53.436 54.937 ;
        RECT 46.628 54.909 53.39 54.983 ;
        RECT 46.582 54.955 53.344 55.029 ;
        RECT 46.536 55.001 53.298 55.075 ;
        RECT 46.49 55.047 53.252 55.121 ;
        RECT 46.444 55.093 53.206 55.167 ;
        RECT 46.398 55.139 53.16 55.213 ;
        RECT 46.352 55.185 53.114 55.259 ;
        RECT 46.306 55.231 53.068 55.305 ;
        RECT 46.26 55.277 53.022 55.351 ;
        RECT 46.214 55.323 52.976 55.397 ;
        RECT 46.168 55.369 52.93 55.443 ;
        RECT 46.122 55.415 52.884 55.489 ;
        RECT 46.076 55.461 52.838 55.535 ;
        RECT 46.03 55.507 52.792 55.581 ;
        RECT 45.984 55.553 52.746 55.627 ;
        RECT 45.938 55.599 52.7 55.673 ;
        RECT 45.892 55.645 52.654 55.719 ;
        RECT 45.846 55.691 52.608 55.765 ;
        RECT 45.8 55.737 52.562 55.811 ;
        RECT 45.754 55.783 52.516 55.857 ;
        RECT 45.708 55.829 52.47 55.903 ;
        RECT 45.662 55.875 52.424 55.949 ;
        RECT 45.616 55.921 52.378 55.995 ;
        RECT 45.57 55.967 52.332 56.041 ;
        RECT 45.524 56.013 52.286 56.087 ;
        RECT 45.478 56.059 52.24 56.133 ;
        RECT 45.432 56.105 52.194 56.179 ;
        RECT 45.386 56.151 52.148 56.225 ;
        RECT 45.34 56.197 52.102 56.271 ;
        RECT 45.294 56.243 52.056 56.317 ;
        RECT 45.248 56.289 52.01 56.363 ;
        RECT 45.202 56.335 51.964 56.409 ;
        RECT 45.156 56.381 51.918 56.455 ;
        RECT 45.11 56.427 51.872 56.501 ;
        RECT 45.064 56.473 51.826 56.547 ;
        RECT 45.018 56.519 51.78 56.593 ;
        RECT 44.972 56.565 51.734 56.639 ;
        RECT 44.926 56.611 51.688 56.685 ;
        RECT 44.88 56.657 51.642 56.731 ;
        RECT 44.834 56.703 51.596 56.777 ;
        RECT 44.788 56.749 51.55 56.823 ;
        RECT 44.742 56.795 51.504 56.869 ;
        RECT 44.696 56.841 51.458 56.915 ;
        RECT 44.65 56.887 51.412 56.961 ;
        RECT 44.604 56.933 51.366 57.007 ;
        RECT 44.558 56.979 51.32 57.053 ;
        RECT 44.512 57.025 51.274 57.099 ;
        RECT 44.466 57.071 51.228 57.145 ;
        RECT 44.42 57.117 51.182 57.191 ;
        RECT 44.374 57.163 51.136 57.237 ;
        RECT 44.328 57.209 51.09 57.283 ;
        RECT 44.282 57.255 51.044 57.329 ;
        RECT 44.236 57.301 50.998 57.375 ;
        RECT 44.19 57.347 50.952 57.421 ;
        RECT 44.144 57.393 50.906 57.467 ;
        RECT 44.098 57.439 50.86 57.513 ;
        RECT 44.052 57.485 50.814 57.559 ;
        RECT 44.006 57.531 50.768 57.605 ;
        RECT 43.96 57.577 50.722 57.651 ;
        RECT 43.914 57.623 50.676 57.697 ;
        RECT 43.868 57.669 50.63 57.743 ;
        RECT 43.822 57.715 50.584 57.789 ;
        RECT 43.776 57.761 50.538 57.835 ;
        RECT 43.73 57.807 50.492 57.881 ;
        RECT 43.684 57.853 50.446 57.927 ;
        RECT 43.638 57.899 50.4 57.973 ;
        RECT 43.592 57.945 50.354 58.019 ;
        RECT 43.546 57.991 50.308 58.065 ;
        RECT 43.5 58.037 50.262 58.111 ;
        RECT 43.454 58.083 50.216 58.157 ;
        RECT 43.408 58.129 50.17 58.203 ;
        RECT 43.362 58.175 50.124 58.249 ;
        RECT 43.316 58.221 50.078 58.295 ;
        RECT 43.27 58.267 50.032 58.341 ;
        RECT 43.224 58.313 49.986 58.387 ;
        RECT 43.178 58.359 49.94 58.433 ;
        RECT 43.132 58.405 49.894 58.479 ;
        RECT 43.086 58.451 49.848 58.525 ;
        RECT 43.04 58.497 49.802 58.571 ;
        RECT 42.994 58.543 49.756 58.617 ;
        RECT 42.948 58.589 49.71 58.663 ;
        RECT 42.902 58.635 49.664 58.709 ;
        RECT 42.856 58.681 49.618 58.755 ;
        RECT 42.81 58.727 49.572 58.801 ;
        RECT 42.764 58.773 49.526 58.847 ;
        RECT 42.718 58.819 49.48 58.893 ;
        RECT 42.672 58.865 49.434 58.939 ;
        RECT 42.626 58.911 49.388 58.985 ;
        RECT 42.58 58.957 49.342 59.031 ;
        RECT 42.534 59.003 49.296 59.077 ;
        RECT 42.488 59.049 49.25 59.123 ;
        RECT 42.442 59.095 49.204 59.169 ;
        RECT 42.396 59.141 49.158 59.215 ;
        RECT 42.35 59.187 49.112 59.261 ;
        RECT 42.304 59.233 49.066 59.307 ;
        RECT 42.258 59.279 49.02 59.353 ;
        RECT 42.212 59.325 48.974 59.399 ;
        RECT 42.166 59.371 48.928 59.445 ;
        RECT 42.12 59.417 48.882 59.491 ;
        RECT 42.074 59.463 48.836 59.537 ;
        RECT 42.028 59.509 48.79 59.583 ;
        RECT 41.982 59.555 48.744 59.629 ;
        RECT 41.936 59.601 48.698 59.675 ;
        RECT 41.89 59.647 48.652 59.721 ;
        RECT 41.844 59.693 48.606 59.767 ;
        RECT 41.798 59.739 48.56 59.813 ;
        RECT 41.752 59.785 48.514 59.859 ;
        RECT 41.706 59.831 48.468 59.905 ;
        RECT 41.66 59.877 48.422 59.951 ;
        RECT 41.614 59.923 48.376 59.997 ;
        RECT 41.568 59.969 48.33 60.043 ;
        RECT 41.522 60.015 48.284 60.089 ;
        RECT 41.476 60.061 48.238 60.135 ;
        RECT 41.43 60.107 48.192 60.181 ;
        RECT 41.384 60.153 48.146 60.227 ;
        RECT 41.338 60.199 48.1 60.273 ;
        RECT 41.292 60.245 48.054 60.319 ;
        RECT 41.246 60.291 48.008 60.365 ;
        RECT 41.184 60.368 47.962 60.411 ;
        RECT 41.2 60.337 47.962 60.411 ;
        RECT 41.138 60.399 47.916 60.457 ;
        RECT 41.092 60.445 47.87 60.503 ;
        RECT 41.046 60.491 47.824 60.549 ;
        RECT 41 60.537 47.778 60.595 ;
        RECT 40.954 60.583 47.732 60.641 ;
        RECT 40.908 60.629 47.686 60.687 ;
        RECT 40.862 60.675 47.64 60.733 ;
        RECT 40.816 60.721 47.594 60.779 ;
        RECT 40.77 60.767 47.548 60.825 ;
        RECT 40.724 60.813 47.502 60.871 ;
        RECT 40.678 60.859 47.456 60.917 ;
        RECT 40.632 60.905 47.41 60.963 ;
        RECT 40.586 60.951 47.364 61.009 ;
        RECT 40.54 60.997 47.318 61.055 ;
        RECT 40.494 61.043 47.272 61.101 ;
        RECT 40.448 61.089 47.226 61.147 ;
        RECT 40.402 61.135 47.18 61.193 ;
        RECT 40.356 61.181 47.134 61.239 ;
        RECT 40.31 61.227 47.088 61.285 ;
        RECT 40.264 61.273 47.042 61.331 ;
        RECT 40.218 61.319 46.996 61.377 ;
        RECT 40.172 61.365 46.95 61.423 ;
        RECT 40.126 61.411 46.904 61.469 ;
        RECT 40.08 61.457 46.858 61.515 ;
        RECT 40.034 61.503 46.812 61.561 ;
        RECT 39.988 61.549 46.766 61.607 ;
        RECT 39.942 61.595 46.72 61.653 ;
        RECT 39.896 61.641 46.674 61.699 ;
        RECT 39.85 61.687 46.628 61.745 ;
        RECT 39.804 61.733 46.582 61.791 ;
        RECT 39.758 61.779 46.536 61.837 ;
        RECT 39.712 61.825 46.49 61.883 ;
        RECT 39.666 61.871 46.444 61.929 ;
        RECT 39.62 61.917 46.398 61.975 ;
        RECT 39.574 61.963 46.352 62.021 ;
        RECT 39.528 62.009 46.306 62.067 ;
        RECT 39.482 62.055 46.26 62.113 ;
        RECT 39.436 62.101 46.214 62.159 ;
        RECT 39.39 62.147 46.168 62.205 ;
        RECT 39.344 62.193 46.122 62.251 ;
        RECT 39.298 62.239 46.076 62.297 ;
        RECT 39.252 62.285 46.03 62.343 ;
        RECT 39.206 62.331 45.984 62.389 ;
        RECT 39.16 62.377 45.938 62.435 ;
        RECT 39.114 62.423 45.892 62.481 ;
        RECT 39.068 62.469 45.846 62.527 ;
        RECT 39.022 62.515 45.8 62.573 ;
        RECT 38.976 62.561 45.754 62.619 ;
        RECT 38.93 62.607 45.708 62.665 ;
        RECT 38.884 62.653 45.662 62.711 ;
        RECT 38.838 62.699 45.616 62.757 ;
        RECT 38.792 62.745 45.57 62.803 ;
        RECT 38.746 62.791 45.524 62.849 ;
        RECT 38.7 62.837 45.478 62.895 ;
        RECT 38.654 62.883 45.432 62.941 ;
        RECT 38.608 62.929 45.386 62.987 ;
        RECT 38.562 62.975 45.34 63.033 ;
        RECT 38.516 63.021 45.294 63.079 ;
        RECT 38.47 63.067 45.248 63.125 ;
        RECT 38.424 63.113 45.202 63.171 ;
        RECT 38.378 63.159 45.156 63.217 ;
        RECT 38.332 63.205 45.11 63.263 ;
        RECT 38.286 63.251 45.064 63.309 ;
        RECT 38.24 63.297 45.018 63.355 ;
        RECT 38.194 63.343 44.972 63.401 ;
        RECT 38.148 63.389 44.926 63.447 ;
        RECT 38.102 63.435 44.88 63.493 ;
        RECT 38.056 63.481 44.834 63.539 ;
        RECT 38.01 63.527 44.788 63.585 ;
        RECT 37.964 63.573 44.742 63.631 ;
        RECT 37.918 63.619 44.696 63.677 ;
        RECT 37.872 63.665 44.65 63.723 ;
        RECT 37.826 63.711 44.604 63.769 ;
        RECT 37.78 63.757 44.558 63.815 ;
        RECT 37.734 63.803 44.512 63.861 ;
        RECT 37.688 63.849 44.466 63.907 ;
        RECT 37.642 63.895 44.42 63.953 ;
        RECT 37.596 63.941 44.374 63.999 ;
        RECT 37.55 63.987 44.328 64.045 ;
        RECT 37.504 64.033 44.282 64.091 ;
        RECT 37.458 64.079 44.236 64.137 ;
        RECT 37.412 64.125 44.19 64.183 ;
        RECT 37.366 64.171 44.144 64.229 ;
        RECT 37.32 64.217 44.098 64.275 ;
        RECT 37.274 64.263 44.052 64.321 ;
        RECT 37.228 64.309 44.006 64.367 ;
        RECT 37.182 64.355 43.96 64.413 ;
        RECT 37.136 64.401 43.914 64.459 ;
        RECT 37.09 64.447 43.868 64.505 ;
        RECT 37.044 64.493 43.822 64.551 ;
        RECT 36.998 64.539 43.776 64.597 ;
        RECT 36.952 64.585 43.73 64.643 ;
        RECT 36.906 64.631 43.684 64.689 ;
        RECT 36.86 64.677 43.638 64.735 ;
        RECT 36.814 64.723 43.592 64.781 ;
        RECT 36.768 64.769 43.546 64.827 ;
        RECT 36.722 64.815 43.5 64.873 ;
        RECT 36.676 64.861 43.454 64.919 ;
        RECT 36.63 64.907 43.408 64.965 ;
        RECT 36.584 64.953 43.362 65.011 ;
        RECT 36.538 64.999 43.316 65.057 ;
        RECT 36.492 65.045 43.27 65.103 ;
        RECT 36.446 65.091 43.224 65.149 ;
        RECT 36.4 65.137 43.178 65.195 ;
        RECT 36.4 65.137 43.132 65.241 ;
        RECT 36.4 65.137 43.086 65.287 ;
        RECT 36.4 65.137 43.04 65.333 ;
        RECT 36.4 65.137 42.994 65.379 ;
        RECT 36.4 65.137 42.948 65.425 ;
        RECT 36.4 65.137 42.902 65.471 ;
        RECT 36.4 65.137 42.856 65.517 ;
        RECT 36.4 65.137 42.81 65.563 ;
        RECT 36.4 65.137 42.764 65.609 ;
        RECT 36.4 65.137 42.718 65.655 ;
        RECT 36.4 65.137 42.672 65.701 ;
        RECT 36.4 65.137 42.626 65.747 ;
        RECT 36.4 65.137 42.58 65.793 ;
        RECT 36.4 65.137 42.534 65.839 ;
        RECT 36.4 65.137 42.488 65.885 ;
        RECT 36.4 65.137 42.442 65.931 ;
        RECT 36.4 65.137 42.396 65.977 ;
        RECT 36.4 65.137 42.35 66.023 ;
        RECT 36.4 65.137 42.304 66.069 ;
        RECT 36.4 65.137 42.258 66.115 ;
        RECT 36.4 65.137 42.212 66.161 ;
        RECT 36.4 65.137 42.166 66.207 ;
        RECT 36.4 65.137 42.12 66.253 ;
        RECT 36.4 65.137 42.074 66.299 ;
        RECT 36.4 65.137 42.028 66.345 ;
        RECT 36.4 65.137 41.982 66.391 ;
        RECT 36.4 65.137 41.936 66.437 ;
        RECT 36.4 65.137 41.89 66.483 ;
        RECT 36.4 65.137 41.844 66.529 ;
        RECT 36.4 65.137 41.798 66.575 ;
        RECT 36.4 65.137 41.752 66.621 ;
        RECT 36.4 65.137 41.706 66.667 ;
        RECT 36.4 65.137 41.66 66.713 ;
        RECT 36.4 65.137 41.614 66.759 ;
        RECT 36.4 65.137 41.568 66.805 ;
        RECT 36.4 65.137 41.522 66.851 ;
        RECT 36.4 65.137 41.476 66.897 ;
        RECT 36.4 65.137 41.43 66.943 ;
        RECT 36.4 65.137 41.384 66.989 ;
        RECT 36.4 65.137 41.338 67.035 ;
        RECT 36.4 65.137 41.292 67.081 ;
        RECT 36.4 65.137 41.246 67.127 ;
        RECT 36.4 65.137 41.2 80 ;
        RECT 60.382 41.155 80 41.2 ;
        RECT 65.16 36.4 80 41.2 ;
        RECT 60.336 41.201 67.15 41.206 ;
        RECT 60.336 41.201 67.138 41.235 ;
        RECT 58.404 43.133 65.16 43.21 ;
        RECT 58.45 43.087 65.206 43.167 ;
        RECT 65.12 36.42 65.16 43.21 ;
        RECT 58.358 43.179 65.12 43.253 ;
        RECT 58.496 43.041 65.252 43.121 ;
        RECT 65.074 36.463 65.12 43.253 ;
        RECT 58.312 43.225 65.074 43.299 ;
        RECT 58.542 42.995 65.298 43.075 ;
        RECT 65.028 36.509 65.074 43.299 ;
        RECT 58.266 43.271 65.028 43.345 ;
        RECT 58.588 42.949 65.344 43.029 ;
        RECT 64.982 36.555 65.028 43.345 ;
        RECT 58.22 43.317 64.982 43.391 ;
        RECT 58.634 42.903 65.39 42.983 ;
        RECT 64.936 36.601 64.982 43.391 ;
        RECT 58.174 43.363 64.936 43.437 ;
        RECT 58.68 42.857 65.436 42.937 ;
        RECT 64.89 36.647 64.936 43.437 ;
        RECT 58.128 43.409 64.89 43.483 ;
        RECT 58.726 42.811 65.482 42.891 ;
        RECT 64.844 36.693 64.89 43.483 ;
        RECT 58.082 43.455 64.844 43.529 ;
        RECT 58.772 42.765 65.528 42.845 ;
        RECT 64.798 36.739 64.844 43.529 ;
        RECT 58.036 43.501 64.798 43.575 ;
        RECT 58.818 42.719 65.574 42.799 ;
        RECT 64.752 36.785 64.798 43.575 ;
        RECT 57.99 43.547 64.752 43.621 ;
        RECT 58.864 42.673 65.62 42.753 ;
        RECT 64.706 36.831 64.752 43.621 ;
        RECT 57.944 43.593 64.706 43.667 ;
        RECT 58.91 42.627 65.666 42.707 ;
        RECT 64.66 36.877 64.706 43.667 ;
        RECT 57.898 43.639 64.66 43.713 ;
        RECT 58.956 42.581 65.712 42.661 ;
        RECT 64.614 36.923 64.66 43.713 ;
        RECT 57.852 43.685 64.614 43.759 ;
        RECT 59.002 42.535 65.758 42.615 ;
        RECT 64.568 36.969 64.614 43.759 ;
        RECT 57.806 43.731 64.568 43.805 ;
        RECT 59.048 42.489 65.804 42.569 ;
        RECT 64.522 37.015 64.568 43.805 ;
        RECT 57.76 43.777 64.522 43.851 ;
        RECT 59.094 42.443 65.85 42.523 ;
        RECT 64.476 37.061 64.522 43.851 ;
        RECT 57.714 43.823 64.476 43.897 ;
        RECT 59.14 42.397 65.896 42.477 ;
        RECT 64.43 37.107 64.476 43.897 ;
        RECT 57.668 43.869 64.43 43.943 ;
        RECT 59.186 42.351 65.942 42.431 ;
        RECT 64.384 37.153 64.43 43.943 ;
        RECT 57.622 43.915 64.384 43.989 ;
        RECT 59.232 42.305 65.988 42.385 ;
        RECT 64.338 37.199 64.384 43.989 ;
        RECT 57.576 43.961 64.338 44.035 ;
        RECT 59.278 42.259 66.034 42.339 ;
        RECT 64.292 37.245 64.338 44.035 ;
        RECT 57.53 44.007 64.292 44.081 ;
        RECT 59.324 42.213 66.08 42.293 ;
        RECT 64.246 37.291 64.292 44.081 ;
        RECT 57.484 44.053 64.246 44.127 ;
        RECT 59.37 42.167 66.126 42.247 ;
        RECT 64.2 37.337 64.246 44.127 ;
        RECT 57.438 44.099 64.2 44.173 ;
        RECT 59.416 42.121 66.172 42.201 ;
        RECT 64.154 37.383 64.2 44.173 ;
        RECT 57.392 44.145 64.154 44.219 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 13.512 51.345 21.884 51.409 ;
        RECT 13.466 51.391 21.838 51.455 ;
        RECT 13.42 51.437 21.792 51.501 ;
        RECT 13.374 51.483 21.746 51.547 ;
        RECT 13.328 51.529 21.7 51.593 ;
        RECT 13.282 51.575 21.654 51.639 ;
        RECT 13.236 51.621 21.608 51.685 ;
        RECT 13.19 51.667 21.562 51.731 ;
        RECT 13.144 51.713 21.516 51.777 ;
        RECT 13.098 51.759 21.47 51.823 ;
        RECT 13.052 51.805 21.424 51.869 ;
        RECT 13.006 51.851 21.378 51.915 ;
        RECT 12.96 51.897 21.332 51.961 ;
        RECT 12.914 51.943 21.286 52.007 ;
        RECT 12.868 51.989 21.24 52.053 ;
        RECT 12.822 52.035 21.194 52.099 ;
        RECT 12.776 52.081 21.148 52.145 ;
        RECT 12.73 52.127 21.102 52.191 ;
        RECT 12.684 52.173 21.056 52.237 ;
        RECT 12.638 52.219 21.01 52.283 ;
        RECT 12.592 52.265 20.964 52.329 ;
        RECT 12.546 52.311 20.918 52.375 ;
        RECT 12.5 52.357 20.872 52.421 ;
        RECT 12.454 52.403 20.826 52.467 ;
        RECT 12.408 52.449 20.78 52.513 ;
        RECT 12.362 52.495 20.734 52.559 ;
        RECT 12.316 52.541 20.688 52.605 ;
        RECT 12.27 52.587 20.642 52.651 ;
        RECT 12.224 52.633 20.596 52.697 ;
        RECT 12.178 52.679 20.55 52.743 ;
        RECT 12.132 52.725 20.504 52.789 ;
        RECT 12.086 52.771 20.458 52.835 ;
        RECT 12.04 52.817 20.412 52.881 ;
        RECT 11.994 52.863 20.366 52.927 ;
        RECT 11.948 52.909 20.32 52.973 ;
        RECT 11.902 52.955 20.274 53.019 ;
        RECT 11.856 53.001 20.228 53.065 ;
        RECT 11.81 53.047 20.182 53.111 ;
        RECT 11.764 53.093 20.136 53.157 ;
        RECT 11.718 53.139 20.09 53.203 ;
        RECT 11.672 53.185 20.044 53.249 ;
        RECT 11.626 53.231 19.998 53.295 ;
        RECT 11.58 53.277 19.952 53.341 ;
        RECT 11.534 53.323 19.906 53.387 ;
        RECT 11.488 53.369 19.86 53.433 ;
        RECT 11.442 53.415 19.814 53.479 ;
        RECT 11.396 53.461 19.768 53.525 ;
        RECT 11.35 53.507 19.722 53.571 ;
        RECT 11.304 53.553 19.676 53.617 ;
        RECT 11.258 53.599 19.63 53.663 ;
        RECT 11.212 53.645 19.584 53.709 ;
        RECT 11.166 53.691 19.538 53.755 ;
        RECT 11.12 53.737 19.492 53.801 ;
        RECT 11.074 53.783 19.446 53.847 ;
        RECT 11.028 53.829 19.4 53.893 ;
        RECT 10.982 53.875 19.354 53.939 ;
        RECT 10.936 53.921 19.308 53.985 ;
        RECT 10.89 53.967 19.262 54.031 ;
        RECT 10.844 54.013 19.216 54.077 ;
        RECT 10.798 54.059 19.17 54.123 ;
        RECT 10.752 54.105 19.124 54.169 ;
        RECT 10.706 54.151 19.078 54.215 ;
        RECT 10.66 54.197 19.032 54.261 ;
        RECT 10.614 54.243 18.986 54.307 ;
        RECT 10.568 54.289 18.94 54.353 ;
        RECT 10.522 54.335 18.894 54.399 ;
        RECT 10.476 54.381 18.848 54.445 ;
        RECT 10.43 54.427 18.802 54.491 ;
        RECT 10.384 54.473 18.756 54.537 ;
        RECT 10.338 54.519 18.71 54.583 ;
        RECT 10.292 54.565 18.664 54.629 ;
        RECT 10.246 54.611 18.618 54.675 ;
        RECT 10.184 54.688 18.572 54.721 ;
        RECT 10.2 54.657 18.572 54.721 ;
        RECT 10.138 54.719 18.526 54.767 ;
        RECT 10.092 54.765 18.48 54.813 ;
        RECT 10.046 54.811 18.434 54.859 ;
        RECT 10 54.857 18.388 54.905 ;
        RECT 9.954 54.903 18.342 54.951 ;
        RECT 9.908 54.949 18.296 54.997 ;
        RECT 9.862 54.995 18.25 55.043 ;
        RECT 9.816 55.041 18.204 55.089 ;
        RECT 9.77 55.087 18.158 55.135 ;
        RECT 9.724 55.133 18.112 55.181 ;
        RECT 9.678 55.179 18.066 55.227 ;
        RECT 9.632 55.225 18.02 55.273 ;
        RECT 9.586 55.271 17.974 55.319 ;
        RECT 9.54 55.317 17.928 55.365 ;
        RECT 9.494 55.363 17.882 55.411 ;
        RECT 9.448 55.409 17.836 55.457 ;
        RECT 9.402 55.455 17.79 55.503 ;
        RECT 9.356 55.501 17.744 55.549 ;
        RECT 9.31 55.547 17.698 55.595 ;
        RECT 9.264 55.593 17.652 55.641 ;
        RECT 9.218 55.639 17.606 55.687 ;
        RECT 9.172 55.685 17.56 55.733 ;
        RECT 9.126 55.731 17.514 55.779 ;
        RECT 9.08 55.777 17.468 55.825 ;
        RECT 9.034 55.823 17.422 55.871 ;
        RECT 8.988 55.869 17.376 55.917 ;
        RECT 8.942 55.915 17.33 55.963 ;
        RECT 8.896 55.961 17.284 56.009 ;
        RECT 8.85 56.007 17.238 56.055 ;
        RECT 8.804 56.053 17.192 56.101 ;
        RECT 8.758 56.099 17.146 56.147 ;
        RECT 8.712 56.145 17.1 56.193 ;
        RECT 8.666 56.191 17.054 56.239 ;
        RECT 8.62 56.237 17.008 56.285 ;
        RECT 8.574 56.283 16.962 56.331 ;
        RECT 8.528 56.329 16.916 56.377 ;
        RECT 8.482 56.375 16.87 56.423 ;
        RECT 8.436 56.421 16.824 56.469 ;
        RECT 8.39 56.467 16.778 56.515 ;
        RECT 8.344 56.513 16.732 56.561 ;
        RECT 8.298 56.559 16.686 56.607 ;
        RECT 8.252 56.605 16.64 56.653 ;
        RECT 8.206 56.651 16.594 56.699 ;
        RECT 8.16 56.697 16.548 56.745 ;
        RECT 8.114 56.743 16.502 56.791 ;
        RECT 8.068 56.789 16.456 56.837 ;
        RECT 8.022 56.835 16.41 56.883 ;
        RECT 7.976 56.881 16.364 56.929 ;
        RECT 7.93 56.927 16.318 56.975 ;
        RECT 7.884 56.973 16.272 57.021 ;
        RECT 7.838 57.019 16.226 57.067 ;
        RECT 7.792 57.065 16.18 57.113 ;
        RECT 7.746 57.111 16.134 57.159 ;
        RECT 7.7 57.157 16.088 57.205 ;
        RECT 7.654 57.203 16.042 57.251 ;
        RECT 7.608 57.249 15.996 57.297 ;
        RECT 7.562 57.295 15.95 57.343 ;
        RECT 7.516 57.341 15.904 57.389 ;
        RECT 7.47 57.387 15.858 57.435 ;
        RECT 7.424 57.433 15.812 57.481 ;
        RECT 7.378 57.479 15.766 57.527 ;
        RECT 7.332 57.525 15.72 57.573 ;
        RECT 7.286 57.571 15.674 57.619 ;
        RECT 7.24 57.617 15.628 57.665 ;
        RECT 7.194 57.663 15.582 57.711 ;
        RECT 7.148 57.709 15.536 57.757 ;
        RECT 7.102 57.755 15.49 57.803 ;
        RECT 7.056 57.801 15.444 57.849 ;
        RECT 7.01 57.847 15.398 57.895 ;
        RECT 6.964 57.893 15.352 57.941 ;
        RECT 6.918 57.939 15.306 57.987 ;
        RECT 6.872 57.985 15.26 58.033 ;
        RECT 6.826 58.031 15.214 58.079 ;
        RECT 6.78 58.077 15.168 58.125 ;
        RECT 6.734 58.123 15.122 58.171 ;
        RECT 6.688 58.169 15.076 58.217 ;
        RECT 6.642 58.215 15.03 58.263 ;
        RECT 6.596 58.261 14.984 58.309 ;
        RECT 6.55 58.307 14.938 58.355 ;
        RECT 6.504 58.353 14.892 58.401 ;
        RECT 6.458 58.399 14.846 58.447 ;
        RECT 6.412 58.445 14.8 58.493 ;
        RECT 6.366 58.491 14.754 58.539 ;
        RECT 6.32 58.537 14.708 58.585 ;
        RECT 6.274 58.583 14.662 58.631 ;
        RECT 6.228 58.629 14.616 58.677 ;
        RECT 6.182 58.675 14.57 58.723 ;
        RECT 6.136 58.721 14.524 58.769 ;
        RECT 6.09 58.767 14.478 58.815 ;
        RECT 6.044 58.813 14.432 58.861 ;
        RECT 5.998 58.859 14.386 58.907 ;
        RECT 5.952 58.905 14.34 58.953 ;
        RECT 5.906 58.951 14.294 58.999 ;
        RECT 5.86 58.997 14.248 59.045 ;
        RECT 5.814 59.043 14.202 59.091 ;
        RECT 5.768 59.089 14.156 59.137 ;
        RECT 5.722 59.135 14.11 59.183 ;
        RECT 5.676 59.181 14.064 59.229 ;
        RECT 5.63 59.227 14.018 59.275 ;
        RECT 5.584 59.273 13.972 59.321 ;
        RECT 5.538 59.319 13.926 59.367 ;
        RECT 5.492 59.365 13.88 59.413 ;
        RECT 5.446 59.411 13.834 59.459 ;
        RECT 5.4 59.457 13.788 59.505 ;
        RECT 5.4 59.457 13.742 59.551 ;
        RECT 5.4 59.457 13.696 59.597 ;
        RECT 5.4 59.457 13.65 59.643 ;
        RECT 5.4 59.457 13.604 59.689 ;
        RECT 5.4 59.457 13.558 59.735 ;
        RECT 5.4 59.457 13.512 59.781 ;
        RECT 5.4 59.457 13.466 59.827 ;
        RECT 5.4 59.457 13.42 59.873 ;
        RECT 5.4 59.457 13.374 59.919 ;
        RECT 5.4 59.457 13.328 59.965 ;
        RECT 5.4 59.457 13.282 60.011 ;
        RECT 5.4 59.457 13.236 60.057 ;
        RECT 5.4 59.457 13.19 60.103 ;
        RECT 5.4 59.457 13.144 60.149 ;
        RECT 5.4 59.457 13.098 60.195 ;
        RECT 5.4 59.457 13.052 60.241 ;
        RECT 5.4 59.457 13.006 60.287 ;
        RECT 5.4 59.457 12.96 60.333 ;
        RECT 5.4 59.457 12.914 60.379 ;
        RECT 5.4 59.457 12.868 60.425 ;
        RECT 5.4 59.457 12.822 60.471 ;
        RECT 5.4 59.457 12.776 60.517 ;
        RECT 5.4 59.457 12.73 60.563 ;
        RECT 5.4 59.457 12.684 60.609 ;
        RECT 5.4 59.457 12.638 60.655 ;
        RECT 5.4 59.457 12.592 60.701 ;
        RECT 5.4 59.457 12.546 60.747 ;
        RECT 5.4 59.457 12.5 60.793 ;
        RECT 5.4 59.457 12.454 60.839 ;
        RECT 5.4 59.457 12.408 60.885 ;
        RECT 5.4 59.457 12.362 60.931 ;
        RECT 5.4 59.457 12.316 60.977 ;
        RECT 5.4 59.457 12.27 61.023 ;
        RECT 5.4 59.457 12.224 61.069 ;
        RECT 5.4 59.457 12.178 61.115 ;
        RECT 5.4 59.457 12.132 61.161 ;
        RECT 5.4 59.457 12.086 61.207 ;
        RECT 5.4 59.457 12.04 61.253 ;
        RECT 5.4 59.457 11.994 61.299 ;
        RECT 5.4 59.457 11.948 61.345 ;
        RECT 5.4 59.457 11.902 61.391 ;
        RECT 5.4 59.457 11.856 61.437 ;
        RECT 5.4 59.457 11.81 61.483 ;
        RECT 5.4 59.457 11.764 61.529 ;
        RECT 5.4 59.457 11.718 61.575 ;
        RECT 5.4 59.457 11.672 61.621 ;
        RECT 5.4 59.457 11.626 61.667 ;
        RECT 5.4 59.457 11.58 61.713 ;
        RECT 5.4 59.457 11.534 61.759 ;
        RECT 5.4 59.457 11.488 61.805 ;
        RECT 5.4 59.457 11.442 61.851 ;
        RECT 5.4 59.457 11.396 61.897 ;
        RECT 5.4 59.457 11.35 61.943 ;
        RECT 5.4 59.457 11.304 61.989 ;
        RECT 5.4 59.457 11.258 62.035 ;
        RECT 5.4 59.457 11.212 62.081 ;
        RECT 5.4 59.457 11.166 62.127 ;
        RECT 5.4 59.457 11.12 62.173 ;
        RECT 5.4 59.457 11.074 62.219 ;
        RECT 5.4 59.457 11.028 62.265 ;
        RECT 5.4 59.457 10.982 62.311 ;
        RECT 5.4 59.457 10.936 62.357 ;
        RECT 5.4 59.457 10.89 62.403 ;
        RECT 5.4 59.457 10.844 62.449 ;
        RECT 5.4 59.457 10.798 62.495 ;
        RECT 5.4 59.457 10.752 62.541 ;
        RECT 5.4 59.457 10.706 62.587 ;
        RECT 5.4 59.457 10.66 62.633 ;
        RECT 5.4 59.457 10.614 62.679 ;
        RECT 5.4 59.457 10.568 62.725 ;
        RECT 5.4 59.457 10.522 62.771 ;
        RECT 5.4 59.457 10.476 62.817 ;
        RECT 5.4 59.457 10.43 62.863 ;
        RECT 5.4 59.457 10.384 62.909 ;
        RECT 5.4 59.457 10.338 62.955 ;
        RECT 5.4 59.457 10.292 63.001 ;
        RECT 5.4 59.457 10.246 63.047 ;
        RECT 5.4 59.457 10.2 80 ;
        RECT 59.48 5.4 80 10.2 ;
        RECT 51.14 13.717 59.526 13.767 ;
        RECT 59.466 5.407 59.48 13.797 ;
        RECT 51.094 13.763 59.466 13.827 ;
        RECT 51.186 13.671 59.572 13.721 ;
        RECT 59.42 5.437 59.466 13.827 ;
        RECT 51.048 13.809 59.42 13.873 ;
        RECT 51.232 13.625 59.618 13.675 ;
        RECT 59.374 5.483 59.42 13.873 ;
        RECT 51.002 13.855 59.374 13.919 ;
        RECT 51.278 13.579 59.664 13.629 ;
        RECT 59.328 5.529 59.374 13.919 ;
        RECT 50.956 13.901 59.328 13.965 ;
        RECT 51.324 13.533 59.71 13.583 ;
        RECT 59.282 5.575 59.328 13.965 ;
        RECT 50.91 13.947 59.282 14.011 ;
        RECT 51.37 13.487 59.756 13.537 ;
        RECT 59.236 5.621 59.282 14.011 ;
        RECT 50.864 13.993 59.236 14.057 ;
        RECT 51.416 13.441 59.802 13.491 ;
        RECT 59.19 5.667 59.236 14.057 ;
        RECT 50.818 14.039 59.19 14.103 ;
        RECT 51.462 13.395 59.848 13.445 ;
        RECT 59.144 5.713 59.19 14.103 ;
        RECT 50.772 14.085 59.144 14.149 ;
        RECT 51.508 13.349 59.894 13.399 ;
        RECT 59.098 5.759 59.144 14.149 ;
        RECT 50.726 14.131 59.098 14.195 ;
        RECT 51.554 13.303 59.94 13.353 ;
        RECT 59.052 5.805 59.098 14.195 ;
        RECT 50.68 14.177 59.052 14.241 ;
        RECT 51.6 13.257 59.986 13.307 ;
        RECT 59.006 5.851 59.052 14.241 ;
        RECT 50.634 14.223 59.006 14.287 ;
        RECT 51.646 13.211 60.032 13.261 ;
        RECT 58.96 5.897 59.006 14.287 ;
        RECT 50.588 14.269 58.96 14.333 ;
        RECT 51.692 13.165 60.078 13.215 ;
        RECT 58.914 5.943 58.96 14.333 ;
        RECT 50.542 14.315 58.914 14.379 ;
        RECT 51.738 13.119 60.124 13.169 ;
        RECT 58.868 5.989 58.914 14.379 ;
        RECT 50.496 14.361 58.868 14.425 ;
        RECT 51.784 13.073 60.17 13.123 ;
        RECT 58.822 6.035 58.868 14.425 ;
        RECT 50.45 14.407 58.822 14.471 ;
        RECT 51.83 13.027 60.216 13.077 ;
        RECT 58.776 6.081 58.822 14.471 ;
        RECT 50.404 14.453 58.776 14.517 ;
        RECT 51.876 12.981 60.262 13.031 ;
        RECT 58.73 6.127 58.776 14.517 ;
        RECT 50.358 14.499 58.73 14.563 ;
        RECT 51.922 12.935 60.308 12.985 ;
        RECT 58.684 6.173 58.73 14.563 ;
        RECT 50.312 14.545 58.684 14.609 ;
        RECT 51.968 12.889 60.354 12.939 ;
        RECT 58.638 6.219 58.684 14.609 ;
        RECT 50.266 14.591 58.638 14.655 ;
        RECT 52.014 12.843 60.4 12.893 ;
        RECT 58.592 6.265 58.638 14.655 ;
        RECT 50.22 14.637 58.592 14.701 ;
        RECT 52.06 12.797 60.446 12.847 ;
        RECT 58.546 6.311 58.592 14.701 ;
        RECT 50.174 14.683 58.546 14.747 ;
        RECT 52.106 12.751 60.492 12.801 ;
        RECT 58.5 6.357 58.546 14.747 ;
        RECT 50.128 14.729 58.5 14.793 ;
        RECT 52.152 12.705 60.538 12.755 ;
        RECT 58.454 6.403 58.5 14.793 ;
        RECT 50.082 14.775 58.454 14.839 ;
        RECT 52.198 12.659 60.584 12.709 ;
        RECT 58.408 6.449 58.454 14.839 ;
        RECT 50.036 14.821 58.408 14.885 ;
        RECT 52.244 12.613 60.63 12.663 ;
        RECT 58.362 6.495 58.408 14.885 ;
        RECT 49.99 14.867 58.362 14.931 ;
        RECT 52.29 12.567 60.676 12.617 ;
        RECT 58.316 6.541 58.362 14.931 ;
        RECT 49.944 14.913 58.316 14.977 ;
        RECT 52.336 12.521 60.722 12.571 ;
        RECT 58.27 6.587 58.316 14.977 ;
        RECT 49.898 14.959 58.27 15.023 ;
        RECT 52.382 12.475 60.768 12.525 ;
        RECT 58.224 6.633 58.27 15.023 ;
        RECT 49.852 15.005 58.224 15.069 ;
        RECT 52.428 12.429 60.814 12.479 ;
        RECT 58.178 6.679 58.224 15.069 ;
        RECT 49.806 15.051 58.178 15.115 ;
        RECT 52.474 12.383 60.86 12.433 ;
        RECT 58.132 6.725 58.178 15.115 ;
        RECT 49.76 15.097 58.132 15.161 ;
        RECT 52.52 12.337 60.906 12.387 ;
        RECT 58.086 6.771 58.132 15.161 ;
        RECT 49.714 15.143 58.086 15.207 ;
        RECT 52.566 12.291 60.952 12.341 ;
        RECT 58.04 6.817 58.086 15.207 ;
        RECT 49.668 15.189 58.04 15.253 ;
        RECT 52.612 12.245 60.998 12.295 ;
        RECT 57.994 6.863 58.04 15.253 ;
        RECT 49.622 15.235 57.994 15.299 ;
        RECT 52.658 12.199 61.044 12.249 ;
        RECT 57.948 6.909 57.994 15.299 ;
        RECT 49.576 15.281 57.948 15.345 ;
        RECT 52.704 12.153 61.09 12.203 ;
        RECT 57.902 6.955 57.948 15.345 ;
        RECT 49.53 15.327 57.902 15.391 ;
        RECT 52.75 12.107 61.136 12.157 ;
        RECT 57.856 7.001 57.902 15.391 ;
        RECT 49.484 15.373 57.856 15.437 ;
        RECT 52.796 12.061 61.182 12.111 ;
        RECT 57.81 7.047 57.856 15.437 ;
        RECT 49.438 15.419 57.81 15.483 ;
        RECT 52.842 12.015 61.228 12.065 ;
        RECT 57.764 7.093 57.81 15.483 ;
        RECT 49.392 15.465 57.764 15.529 ;
        RECT 52.888 11.969 61.274 12.019 ;
        RECT 57.718 7.139 57.764 15.529 ;
        RECT 49.346 15.511 57.718 15.575 ;
        RECT 52.934 11.923 61.32 11.973 ;
        RECT 57.672 7.185 57.718 15.575 ;
        RECT 49.3 15.557 57.672 15.621 ;
        RECT 52.98 11.877 61.366 11.927 ;
        RECT 57.626 7.231 57.672 15.621 ;
        RECT 49.254 15.603 57.626 15.667 ;
        RECT 53.026 11.831 61.412 11.881 ;
        RECT 57.58 7.277 57.626 15.667 ;
        RECT 49.208 15.649 57.58 15.713 ;
        RECT 53.072 11.785 61.458 11.835 ;
        RECT 57.534 7.323 57.58 15.713 ;
        RECT 49.162 15.695 57.534 15.759 ;
        RECT 53.118 11.739 61.504 11.789 ;
        RECT 57.488 7.369 57.534 15.759 ;
        RECT 49.116 15.741 57.488 15.805 ;
        RECT 53.164 11.693 61.55 11.743 ;
        RECT 57.442 7.415 57.488 15.805 ;
        RECT 49.07 15.787 57.442 15.851 ;
        RECT 53.21 11.647 61.596 11.697 ;
        RECT 57.396 7.461 57.442 15.851 ;
        RECT 49.024 15.833 57.396 15.897 ;
        RECT 53.256 11.601 61.642 11.651 ;
        RECT 57.35 7.507 57.396 15.897 ;
        RECT 48.978 15.879 57.35 15.943 ;
        RECT 53.302 11.555 61.688 11.605 ;
        RECT 57.304 7.553 57.35 15.943 ;
        RECT 48.932 15.925 57.304 15.989 ;
        RECT 53.348 11.509 61.734 11.559 ;
        RECT 57.258 7.599 57.304 15.989 ;
        RECT 48.886 15.971 57.258 16.035 ;
        RECT 53.394 11.463 61.78 11.513 ;
        RECT 57.212 7.645 57.258 16.035 ;
        RECT 48.84 16.017 57.212 16.081 ;
        RECT 53.44 11.417 61.826 11.467 ;
        RECT 57.166 7.691 57.212 16.081 ;
        RECT 48.794 16.063 57.166 16.127 ;
        RECT 53.486 11.371 61.872 11.421 ;
        RECT 57.12 7.737 57.166 16.127 ;
        RECT 48.748 16.109 57.12 16.173 ;
        RECT 53.532 11.325 61.918 11.375 ;
        RECT 57.074 7.783 57.12 16.173 ;
        RECT 48.702 16.155 57.074 16.219 ;
        RECT 53.578 11.279 61.964 11.329 ;
        RECT 57.028 7.829 57.074 16.219 ;
        RECT 48.656 16.201 57.028 16.265 ;
        RECT 53.624 11.233 62.01 11.283 ;
        RECT 56.982 7.875 57.028 16.265 ;
        RECT 48.61 16.247 56.982 16.311 ;
        RECT 53.67 11.187 62.056 11.237 ;
        RECT 56.936 7.921 56.982 16.311 ;
        RECT 48.564 16.293 56.936 16.357 ;
        RECT 53.716 11.141 62.102 11.191 ;
        RECT 56.89 7.967 56.936 16.357 ;
        RECT 48.518 16.339 56.89 16.403 ;
        RECT 53.762 11.095 62.148 11.145 ;
        RECT 56.844 8.013 56.89 16.403 ;
        RECT 48.472 16.385 56.844 16.449 ;
        RECT 53.808 11.049 62.194 11.099 ;
        RECT 56.798 8.059 56.844 16.449 ;
        RECT 48.426 16.431 56.798 16.495 ;
        RECT 53.854 11.003 62.24 11.053 ;
        RECT 56.752 8.105 56.798 16.495 ;
        RECT 48.38 16.477 56.752 16.541 ;
        RECT 53.9 10.957 62.286 11.007 ;
        RECT 56.706 8.151 56.752 16.541 ;
        RECT 48.334 16.523 56.706 16.587 ;
        RECT 53.946 10.911 62.332 10.961 ;
        RECT 56.66 8.197 56.706 16.587 ;
        RECT 48.288 16.569 56.66 16.633 ;
        RECT 53.992 10.865 62.378 10.915 ;
        RECT 56.614 8.243 56.66 16.633 ;
        RECT 48.242 16.615 56.614 16.679 ;
        RECT 54.038 10.819 62.424 10.869 ;
        RECT 56.568 8.289 56.614 16.679 ;
        RECT 48.196 16.661 56.568 16.725 ;
        RECT 54.084 10.773 62.47 10.823 ;
        RECT 56.522 8.335 56.568 16.725 ;
        RECT 48.15 16.707 56.522 16.771 ;
        RECT 54.13 10.727 62.516 10.777 ;
        RECT 56.476 8.381 56.522 16.771 ;
        RECT 48.104 16.753 56.476 16.817 ;
        RECT 54.176 10.681 62.562 10.731 ;
        RECT 56.43 8.427 56.476 16.817 ;
        RECT 48.058 16.799 56.43 16.863 ;
        RECT 54.222 10.635 62.608 10.685 ;
        RECT 56.384 8.473 56.43 16.863 ;
        RECT 48.012 16.845 56.384 16.909 ;
        RECT 54.268 10.589 62.654 10.639 ;
        RECT 56.338 8.519 56.384 16.909 ;
        RECT 47.966 16.891 56.338 16.955 ;
        RECT 54.314 10.543 62.7 10.593 ;
        RECT 56.292 8.565 56.338 16.955 ;
        RECT 47.92 16.937 56.292 17.001 ;
        RECT 54.36 10.497 62.746 10.547 ;
        RECT 56.246 8.611 56.292 17.001 ;
        RECT 47.874 16.983 56.246 17.047 ;
        RECT 54.406 10.451 62.792 10.501 ;
        RECT 56.2 8.657 56.246 17.047 ;
        RECT 47.828 17.029 56.2 17.093 ;
        RECT 54.452 10.405 62.838 10.455 ;
        RECT 56.154 8.703 56.2 17.093 ;
        RECT 47.782 17.075 56.154 17.139 ;
        RECT 54.498 10.359 62.884 10.409 ;
        RECT 56.108 8.749 56.154 17.139 ;
        RECT 47.736 17.121 56.108 17.185 ;
        RECT 54.544 10.313 62.93 10.363 ;
        RECT 56.062 8.795 56.108 17.185 ;
        RECT 47.69 17.167 56.062 17.231 ;
        RECT 54.59 10.267 62.976 10.317 ;
        RECT 56.016 8.841 56.062 17.231 ;
        RECT 47.644 17.213 56.016 17.277 ;
        RECT 54.636 10.221 63.022 10.271 ;
        RECT 55.97 8.887 56.016 17.277 ;
        RECT 47.598 17.259 55.97 17.323 ;
        RECT 54.682 10.175 63.068 10.224 ;
        RECT 55.924 8.933 55.97 17.323 ;
        RECT 47.552 17.305 55.924 17.369 ;
        RECT 54.728 10.129 80 10.2 ;
        RECT 55.878 8.979 55.924 17.369 ;
        RECT 47.506 17.351 55.878 17.415 ;
        RECT 54.774 10.083 80 10.2 ;
        RECT 55.832 9.025 55.878 17.415 ;
        RECT 47.46 17.397 55.832 17.461 ;
        RECT 54.82 10.037 80 10.2 ;
        RECT 55.786 9.071 55.832 17.461 ;
        RECT 47.414 17.443 55.786 17.507 ;
        RECT 54.866 9.991 80 10.2 ;
        RECT 55.74 9.117 55.786 17.507 ;
        RECT 47.368 17.489 55.74 17.553 ;
        RECT 54.912 9.945 80 10.2 ;
        RECT 55.694 9.163 55.74 17.553 ;
        RECT 47.322 17.535 55.694 17.599 ;
        RECT 54.958 9.899 80 10.2 ;
        RECT 55.648 9.209 55.694 17.599 ;
        RECT 47.276 17.581 55.648 17.645 ;
        RECT 55.004 9.853 80 10.2 ;
        RECT 55.602 9.255 55.648 17.645 ;
        RECT 47.23 17.627 55.602 17.691 ;
        RECT 55.05 9.807 80 10.2 ;
        RECT 55.556 9.301 55.602 17.691 ;
        RECT 47.184 17.673 55.556 17.737 ;
        RECT 55.096 9.761 80 10.2 ;
        RECT 55.51 9.347 55.556 17.737 ;
        RECT 47.138 17.719 55.51 17.783 ;
        RECT 55.142 9.715 80 10.2 ;
        RECT 55.464 9.393 55.51 17.783 ;
        RECT 47.092 17.765 55.464 17.829 ;
        RECT 55.188 9.669 80 10.2 ;
        RECT 55.418 9.439 55.464 17.829 ;
        RECT 47.046 17.811 55.418 17.875 ;
        RECT 55.234 9.623 80 10.2 ;
        RECT 55.372 9.485 55.418 17.875 ;
        RECT 47 17.857 55.372 17.921 ;
        RECT 55.28 9.577 80 10.2 ;
        RECT 55.326 9.531 55.372 17.921 ;
        RECT 46.954 17.903 55.326 17.967 ;
        RECT 46.908 17.949 55.28 18.013 ;
        RECT 46.862 17.995 55.234 18.059 ;
        RECT 46.816 18.041 55.188 18.105 ;
        RECT 46.77 18.087 55.142 18.151 ;
        RECT 46.724 18.133 55.096 18.197 ;
        RECT 46.678 18.179 55.05 18.243 ;
        RECT 46.632 18.225 55.004 18.289 ;
        RECT 46.586 18.271 54.958 18.335 ;
        RECT 46.54 18.317 54.912 18.381 ;
        RECT 46.494 18.363 54.866 18.427 ;
        RECT 46.448 18.409 54.82 18.473 ;
        RECT 46.402 18.455 54.774 18.519 ;
        RECT 46.356 18.501 54.728 18.565 ;
        RECT 46.31 18.547 54.682 18.611 ;
        RECT 46.264 18.593 54.636 18.657 ;
        RECT 46.218 18.639 54.59 18.703 ;
        RECT 46.172 18.685 54.544 18.749 ;
        RECT 46.126 18.731 54.498 18.795 ;
        RECT 46.08 18.777 54.452 18.841 ;
        RECT 46.034 18.823 54.406 18.887 ;
        RECT 45.988 18.869 54.36 18.933 ;
        RECT 45.942 18.915 54.314 18.979 ;
        RECT 45.896 18.961 54.268 19.025 ;
        RECT 45.85 19.007 54.222 19.071 ;
        RECT 45.804 19.053 54.176 19.117 ;
        RECT 45.758 19.099 54.13 19.163 ;
        RECT 45.712 19.145 54.084 19.209 ;
        RECT 45.666 19.191 54.038 19.255 ;
        RECT 45.62 19.237 53.992 19.301 ;
        RECT 45.574 19.283 53.946 19.347 ;
        RECT 45.528 19.329 53.9 19.393 ;
        RECT 45.482 19.375 53.854 19.439 ;
        RECT 45.436 19.421 53.808 19.485 ;
        RECT 45.39 19.467 53.762 19.531 ;
        RECT 45.344 19.513 53.716 19.577 ;
        RECT 45.298 19.559 53.67 19.623 ;
        RECT 45.252 19.605 53.624 19.669 ;
        RECT 45.206 19.651 53.578 19.715 ;
        RECT 45.16 19.697 53.532 19.761 ;
        RECT 45.114 19.743 53.486 19.807 ;
        RECT 45.068 19.789 53.44 19.853 ;
        RECT 45.022 19.835 53.394 19.899 ;
        RECT 44.976 19.881 53.348 19.945 ;
        RECT 44.93 19.927 53.302 19.991 ;
        RECT 44.884 19.973 53.256 20.037 ;
        RECT 44.838 20.019 53.21 20.083 ;
        RECT 44.792 20.065 53.164 20.129 ;
        RECT 44.746 20.111 53.118 20.175 ;
        RECT 44.7 20.157 53.072 20.221 ;
        RECT 44.654 20.203 53.026 20.267 ;
        RECT 44.608 20.249 52.98 20.313 ;
        RECT 44.562 20.295 52.934 20.359 ;
        RECT 44.516 20.341 52.888 20.405 ;
        RECT 44.47 20.387 52.842 20.451 ;
        RECT 44.424 20.433 52.796 20.497 ;
        RECT 44.378 20.479 52.75 20.543 ;
        RECT 44.332 20.525 52.704 20.589 ;
        RECT 44.286 20.571 52.658 20.635 ;
        RECT 44.24 20.617 52.612 20.681 ;
        RECT 44.194 20.663 52.566 20.727 ;
        RECT 44.148 20.709 52.52 20.773 ;
        RECT 44.102 20.755 52.474 20.819 ;
        RECT 44.056 20.801 52.428 20.865 ;
        RECT 44.01 20.847 52.382 20.911 ;
        RECT 43.964 20.893 52.336 20.957 ;
        RECT 43.918 20.939 52.29 21.003 ;
        RECT 43.872 20.985 52.244 21.049 ;
        RECT 43.826 21.031 52.198 21.095 ;
        RECT 43.78 21.077 52.152 21.141 ;
        RECT 43.734 21.123 52.106 21.187 ;
        RECT 43.688 21.169 52.06 21.233 ;
        RECT 43.642 21.215 52.014 21.279 ;
        RECT 43.596 21.261 51.968 21.325 ;
        RECT 43.55 21.307 51.922 21.371 ;
        RECT 43.504 21.353 51.876 21.417 ;
        RECT 43.458 21.399 51.83 21.463 ;
        RECT 43.412 21.445 51.784 21.509 ;
        RECT 43.366 21.491 51.738 21.555 ;
        RECT 43.32 21.537 51.692 21.601 ;
        RECT 43.274 21.583 51.646 21.647 ;
        RECT 43.228 21.629 51.6 21.693 ;
        RECT 43.182 21.675 51.554 21.739 ;
        RECT 43.136 21.721 51.508 21.785 ;
        RECT 43.09 21.767 51.462 21.831 ;
        RECT 43.044 21.813 51.416 21.877 ;
        RECT 42.998 21.859 51.37 21.923 ;
        RECT 42.952 21.905 51.324 21.969 ;
        RECT 42.906 21.951 51.278 22.015 ;
        RECT 42.86 21.997 51.232 22.061 ;
        RECT 42.814 22.043 51.186 22.107 ;
        RECT 42.768 22.089 51.14 22.153 ;
        RECT 42.722 22.135 51.094 22.199 ;
        RECT 42.676 22.181 51.048 22.245 ;
        RECT 42.63 22.227 51.002 22.291 ;
        RECT 42.584 22.273 50.956 22.337 ;
        RECT 42.538 22.319 50.91 22.383 ;
        RECT 42.492 22.365 50.864 22.429 ;
        RECT 42.446 22.411 50.818 22.475 ;
        RECT 42.4 22.457 50.772 22.521 ;
        RECT 42.354 22.503 50.726 22.567 ;
        RECT 42.308 22.549 50.68 22.613 ;
        RECT 42.262 22.595 50.634 22.659 ;
        RECT 42.216 22.641 50.588 22.705 ;
        RECT 42.17 22.687 50.542 22.751 ;
        RECT 42.124 22.733 50.496 22.797 ;
        RECT 42.078 22.779 50.45 22.843 ;
        RECT 42.032 22.825 50.404 22.889 ;
        RECT 41.986 22.871 50.358 22.935 ;
        RECT 41.94 22.917 50.312 22.981 ;
        RECT 41.894 22.963 50.266 23.027 ;
        RECT 41.848 23.009 50.22 23.073 ;
        RECT 41.802 23.055 50.174 23.119 ;
        RECT 41.756 23.101 50.128 23.165 ;
        RECT 41.71 23.147 50.082 23.211 ;
        RECT 41.664 23.193 50.036 23.257 ;
        RECT 41.618 23.239 49.99 23.303 ;
        RECT 41.572 23.285 49.944 23.349 ;
        RECT 41.526 23.331 49.898 23.395 ;
        RECT 41.48 23.377 49.852 23.441 ;
        RECT 41.434 23.423 49.806 23.487 ;
        RECT 41.388 23.469 49.76 23.533 ;
        RECT 41.342 23.515 49.714 23.579 ;
        RECT 41.296 23.561 49.668 23.625 ;
        RECT 41.25 23.607 49.622 23.671 ;
        RECT 41.204 23.653 49.576 23.717 ;
        RECT 41.158 23.699 49.53 23.763 ;
        RECT 41.112 23.745 49.484 23.809 ;
        RECT 41.066 23.791 49.438 23.855 ;
        RECT 41.02 23.837 49.392 23.901 ;
        RECT 40.974 23.883 49.346 23.947 ;
        RECT 40.928 23.929 49.3 23.993 ;
        RECT 40.882 23.975 49.254 24.039 ;
        RECT 40.836 24.021 49.208 24.085 ;
        RECT 40.79 24.067 49.162 24.131 ;
        RECT 40.744 24.113 49.116 24.177 ;
        RECT 40.698 24.159 49.07 24.223 ;
        RECT 40.652 24.205 49.024 24.269 ;
        RECT 40.606 24.251 48.978 24.315 ;
        RECT 40.56 24.297 48.932 24.361 ;
        RECT 40.514 24.343 48.886 24.407 ;
        RECT 40.468 24.389 48.84 24.453 ;
        RECT 40.422 24.435 48.794 24.499 ;
        RECT 40.376 24.481 48.748 24.545 ;
        RECT 40.33 24.527 48.702 24.591 ;
        RECT 40.284 24.573 48.656 24.637 ;
        RECT 40.238 24.619 48.61 24.683 ;
        RECT 40.192 24.665 48.564 24.729 ;
        RECT 40.146 24.711 48.518 24.775 ;
        RECT 40.1 24.757 48.472 24.821 ;
        RECT 40.054 24.803 48.426 24.867 ;
        RECT 40.008 24.849 48.38 24.913 ;
        RECT 39.962 24.895 48.334 24.959 ;
        RECT 39.916 24.941 48.288 25.005 ;
        RECT 39.87 24.987 48.242 25.051 ;
        RECT 39.824 25.033 48.196 25.097 ;
        RECT 39.778 25.079 48.15 25.143 ;
        RECT 39.732 25.125 48.104 25.189 ;
        RECT 39.686 25.171 48.058 25.235 ;
        RECT 39.64 25.217 48.012 25.281 ;
        RECT 39.594 25.263 47.966 25.327 ;
        RECT 39.548 25.309 47.92 25.373 ;
        RECT 39.502 25.355 47.874 25.419 ;
        RECT 39.456 25.401 47.828 25.465 ;
        RECT 39.41 25.447 47.782 25.511 ;
        RECT 39.364 25.493 47.736 25.557 ;
        RECT 39.318 25.539 47.69 25.603 ;
        RECT 39.272 25.585 47.644 25.649 ;
        RECT 39.226 25.631 47.598 25.695 ;
        RECT 39.18 25.677 47.552 25.741 ;
        RECT 39.134 25.723 47.506 25.787 ;
        RECT 39.088 25.769 47.46 25.833 ;
        RECT 39.042 25.815 47.414 25.879 ;
        RECT 38.996 25.861 47.368 25.925 ;
        RECT 38.95 25.907 47.322 25.971 ;
        RECT 38.904 25.953 47.276 26.017 ;
        RECT 38.858 25.999 47.23 26.063 ;
        RECT 38.812 26.045 47.184 26.109 ;
        RECT 38.766 26.091 47.138 26.155 ;
        RECT 38.72 26.137 47.092 26.201 ;
        RECT 38.674 26.183 47.046 26.247 ;
        RECT 38.628 26.229 47 26.293 ;
        RECT 38.582 26.275 46.954 26.339 ;
        RECT 38.536 26.321 46.908 26.385 ;
        RECT 38.49 26.367 46.862 26.431 ;
        RECT 38.444 26.413 46.816 26.477 ;
        RECT 38.398 26.459 46.77 26.523 ;
        RECT 38.352 26.505 46.724 26.569 ;
        RECT 38.306 26.551 46.678 26.615 ;
        RECT 38.26 26.597 46.632 26.661 ;
        RECT 38.214 26.643 46.586 26.707 ;
        RECT 38.168 26.689 46.54 26.753 ;
        RECT 38.122 26.735 46.494 26.799 ;
        RECT 38.076 26.781 46.448 26.845 ;
        RECT 38.03 26.827 46.402 26.891 ;
        RECT 37.984 26.873 46.356 26.937 ;
        RECT 37.938 26.919 46.31 26.983 ;
        RECT 37.892 26.965 46.264 27.029 ;
        RECT 37.846 27.011 46.218 27.075 ;
        RECT 37.8 27.057 46.172 27.121 ;
        RECT 37.754 27.103 46.126 27.167 ;
        RECT 37.708 27.149 46.08 27.213 ;
        RECT 37.662 27.195 46.034 27.259 ;
        RECT 37.616 27.241 45.988 27.305 ;
        RECT 37.57 27.287 45.942 27.351 ;
        RECT 37.524 27.333 45.896 27.397 ;
        RECT 37.478 27.379 45.85 27.443 ;
        RECT 37.432 27.425 45.804 27.489 ;
        RECT 37.386 27.471 45.758 27.535 ;
        RECT 37.34 27.517 45.712 27.581 ;
        RECT 37.294 27.563 45.666 27.627 ;
        RECT 37.248 27.609 45.62 27.673 ;
        RECT 37.202 27.655 45.574 27.719 ;
        RECT 37.156 27.701 45.528 27.765 ;
        RECT 37.11 27.747 45.482 27.811 ;
        RECT 37.064 27.793 45.436 27.857 ;
        RECT 37.018 27.839 45.39 27.903 ;
        RECT 36.972 27.885 45.344 27.949 ;
        RECT 36.926 27.931 45.298 27.995 ;
        RECT 36.88 27.977 45.252 28.041 ;
        RECT 36.834 28.023 45.206 28.087 ;
        RECT 36.788 28.069 45.16 28.133 ;
        RECT 36.742 28.115 45.114 28.179 ;
        RECT 36.696 28.161 45.068 28.225 ;
        RECT 36.65 28.207 45.022 28.271 ;
        RECT 36.604 28.253 44.976 28.317 ;
        RECT 36.558 28.299 44.93 28.363 ;
        RECT 36.512 28.345 44.884 28.409 ;
        RECT 36.466 28.391 44.838 28.455 ;
        RECT 36.42 28.437 44.792 28.501 ;
        RECT 36.374 28.483 44.746 28.547 ;
        RECT 36.328 28.529 44.7 28.593 ;
        RECT 36.282 28.575 44.654 28.639 ;
        RECT 36.236 28.621 44.608 28.685 ;
        RECT 36.19 28.667 44.562 28.731 ;
        RECT 36.144 28.713 44.516 28.777 ;
        RECT 36.098 28.759 44.47 28.823 ;
        RECT 36.052 28.805 44.424 28.869 ;
        RECT 36.006 28.851 44.378 28.915 ;
        RECT 35.96 28.897 44.332 28.961 ;
        RECT 35.914 28.943 44.286 29.007 ;
        RECT 35.868 28.989 44.24 29.053 ;
        RECT 35.822 29.035 44.194 29.099 ;
        RECT 35.776 29.081 44.148 29.145 ;
        RECT 35.73 29.127 44.102 29.191 ;
        RECT 35.684 29.173 44.056 29.237 ;
        RECT 35.638 29.219 44.01 29.283 ;
        RECT 35.592 29.265 43.964 29.329 ;
        RECT 35.546 29.311 43.918 29.375 ;
        RECT 35.5 29.357 43.872 29.421 ;
        RECT 35.454 29.403 43.826 29.467 ;
        RECT 35.408 29.449 43.78 29.513 ;
        RECT 35.362 29.495 43.734 29.559 ;
        RECT 35.316 29.541 43.688 29.605 ;
        RECT 35.27 29.587 43.642 29.651 ;
        RECT 35.224 29.633 43.596 29.697 ;
        RECT 35.178 29.679 43.55 29.743 ;
        RECT 35.132 29.725 43.504 29.789 ;
        RECT 35.086 29.771 43.458 29.835 ;
        RECT 35.04 29.817 43.412 29.881 ;
        RECT 34.994 29.863 43.366 29.927 ;
        RECT 34.948 29.909 43.32 29.973 ;
        RECT 34.902 29.955 43.274 30.019 ;
        RECT 34.856 30.001 43.228 30.065 ;
        RECT 34.81 30.047 43.182 30.111 ;
        RECT 34.764 30.093 43.136 30.157 ;
        RECT 34.718 30.139 43.09 30.203 ;
        RECT 34.672 30.185 43.044 30.249 ;
        RECT 34.626 30.231 42.998 30.295 ;
        RECT 34.58 30.277 42.952 30.341 ;
        RECT 34.534 30.323 42.906 30.387 ;
        RECT 34.488 30.369 42.86 30.433 ;
        RECT 34.442 30.415 42.814 30.479 ;
        RECT 34.396 30.461 42.768 30.525 ;
        RECT 34.35 30.507 42.722 30.571 ;
        RECT 34.304 30.553 42.676 30.617 ;
        RECT 34.258 30.599 42.63 30.663 ;
        RECT 34.212 30.645 42.584 30.709 ;
        RECT 34.166 30.691 42.538 30.755 ;
        RECT 34.12 30.737 42.492 30.801 ;
        RECT 34.074 30.783 42.446 30.847 ;
        RECT 34.028 30.829 42.4 30.893 ;
        RECT 33.982 30.875 42.354 30.939 ;
        RECT 33.936 30.921 42.308 30.985 ;
        RECT 33.89 30.967 42.262 31.031 ;
        RECT 33.844 31.013 42.216 31.077 ;
        RECT 33.798 31.059 42.17 31.123 ;
        RECT 33.752 31.105 42.124 31.169 ;
        RECT 33.706 31.151 42.078 31.215 ;
        RECT 33.66 31.197 42.032 31.261 ;
        RECT 33.614 31.243 41.986 31.307 ;
        RECT 33.568 31.289 41.94 31.353 ;
        RECT 33.522 31.335 41.894 31.399 ;
        RECT 33.476 31.381 41.848 31.445 ;
        RECT 33.43 31.427 41.802 31.491 ;
        RECT 33.384 31.473 41.756 31.537 ;
        RECT 33.338 31.519 41.71 31.583 ;
        RECT 33.292 31.565 41.664 31.629 ;
        RECT 33.246 31.611 41.618 31.675 ;
        RECT 33.2 31.657 41.572 31.721 ;
        RECT 33.154 31.703 41.526 31.767 ;
        RECT 33.108 31.749 41.48 31.813 ;
        RECT 33.062 31.795 41.434 31.859 ;
        RECT 33.016 31.841 41.388 31.905 ;
        RECT 32.97 31.887 41.342 31.951 ;
        RECT 32.924 31.933 41.296 31.997 ;
        RECT 32.878 31.979 41.25 32.043 ;
        RECT 32.832 32.025 41.204 32.089 ;
        RECT 32.786 32.071 41.158 32.135 ;
        RECT 32.74 32.117 41.112 32.181 ;
        RECT 32.694 32.163 41.066 32.227 ;
        RECT 32.648 32.209 41.02 32.273 ;
        RECT 32.602 32.255 40.974 32.319 ;
        RECT 32.556 32.301 40.928 32.365 ;
        RECT 32.51 32.347 40.882 32.411 ;
        RECT 32.464 32.393 40.836 32.457 ;
        RECT 32.418 32.439 40.79 32.503 ;
        RECT 32.372 32.485 40.744 32.549 ;
        RECT 32.326 32.531 40.698 32.595 ;
        RECT 32.28 32.577 40.652 32.641 ;
        RECT 32.234 32.623 40.606 32.687 ;
        RECT 32.188 32.669 40.56 32.733 ;
        RECT 32.142 32.715 40.514 32.779 ;
        RECT 32.096 32.761 40.468 32.825 ;
        RECT 32.05 32.807 40.422 32.871 ;
        RECT 32.004 32.853 40.376 32.917 ;
        RECT 31.958 32.899 40.33 32.963 ;
        RECT 31.912 32.945 40.284 33.009 ;
        RECT 31.866 32.991 40.238 33.055 ;
        RECT 31.82 33.037 40.192 33.101 ;
        RECT 31.774 33.083 40.146 33.147 ;
        RECT 31.728 33.129 40.1 33.193 ;
        RECT 31.682 33.175 40.054 33.239 ;
        RECT 31.636 33.221 40.008 33.285 ;
        RECT 31.59 33.267 39.962 33.331 ;
        RECT 31.544 33.313 39.916 33.377 ;
        RECT 31.498 33.359 39.87 33.423 ;
        RECT 31.452 33.405 39.824 33.469 ;
        RECT 31.406 33.451 39.778 33.515 ;
        RECT 31.36 33.497 39.732 33.561 ;
        RECT 31.314 33.543 39.686 33.607 ;
        RECT 31.268 33.589 39.64 33.653 ;
        RECT 31.222 33.635 39.594 33.699 ;
        RECT 31.176 33.681 39.548 33.745 ;
        RECT 31.13 33.727 39.502 33.791 ;
        RECT 31.084 33.773 39.456 33.837 ;
        RECT 31.038 33.819 39.41 33.883 ;
        RECT 30.992 33.865 39.364 33.929 ;
        RECT 30.946 33.911 39.318 33.975 ;
        RECT 30.9 33.957 39.272 34.021 ;
        RECT 30.854 34.003 39.226 34.067 ;
        RECT 30.808 34.049 39.18 34.113 ;
        RECT 30.762 34.095 39.134 34.159 ;
        RECT 30.716 34.141 39.088 34.205 ;
        RECT 30.67 34.187 39.042 34.251 ;
        RECT 30.624 34.233 38.996 34.297 ;
        RECT 30.578 34.279 38.95 34.343 ;
        RECT 30.532 34.325 38.904 34.389 ;
        RECT 30.486 34.371 38.858 34.435 ;
        RECT 30.44 34.417 38.812 34.481 ;
        RECT 30.394 34.463 38.766 34.527 ;
        RECT 30.348 34.509 38.72 34.573 ;
        RECT 30.302 34.555 38.674 34.619 ;
        RECT 30.256 34.601 38.628 34.665 ;
        RECT 30.21 34.647 38.582 34.711 ;
        RECT 30.164 34.693 38.536 34.757 ;
        RECT 30.118 34.739 38.49 34.803 ;
        RECT 30.072 34.785 38.444 34.849 ;
        RECT 30.026 34.831 38.398 34.895 ;
        RECT 29.98 34.877 38.352 34.941 ;
        RECT 29.934 34.923 38.306 34.987 ;
        RECT 29.888 34.969 38.26 35.033 ;
        RECT 29.842 35.015 38.214 35.079 ;
        RECT 29.796 35.061 38.168 35.125 ;
        RECT 29.75 35.107 38.122 35.171 ;
        RECT 29.704 35.153 38.076 35.217 ;
        RECT 29.658 35.199 38.03 35.263 ;
        RECT 29.612 35.245 37.984 35.309 ;
        RECT 29.566 35.291 37.938 35.355 ;
        RECT 29.52 35.337 37.892 35.401 ;
        RECT 29.474 35.383 37.846 35.447 ;
        RECT 29.428 35.429 37.8 35.493 ;
        RECT 29.382 35.475 37.754 35.539 ;
        RECT 29.336 35.521 37.708 35.585 ;
        RECT 29.29 35.567 37.662 35.631 ;
        RECT 29.244 35.613 37.616 35.677 ;
        RECT 29.198 35.659 37.57 35.723 ;
        RECT 29.152 35.705 37.524 35.769 ;
        RECT 29.106 35.751 37.478 35.815 ;
        RECT 29.06 35.797 37.432 35.861 ;
        RECT 29.014 35.843 37.386 35.907 ;
        RECT 28.968 35.889 37.34 35.953 ;
        RECT 28.922 35.935 37.294 35.999 ;
        RECT 28.876 35.981 37.248 36.045 ;
        RECT 28.83 36.027 37.202 36.091 ;
        RECT 28.784 36.073 37.156 36.137 ;
        RECT 28.738 36.119 37.11 36.183 ;
        RECT 28.692 36.165 37.064 36.229 ;
        RECT 28.646 36.211 37.018 36.275 ;
        RECT 28.6 36.257 36.972 36.321 ;
        RECT 28.554 36.303 36.926 36.367 ;
        RECT 28.508 36.349 36.88 36.413 ;
        RECT 28.462 36.395 36.834 36.459 ;
        RECT 28.416 36.441 36.788 36.505 ;
        RECT 28.37 36.487 36.742 36.551 ;
        RECT 28.324 36.533 36.696 36.597 ;
        RECT 28.278 36.579 36.65 36.643 ;
        RECT 28.232 36.625 36.604 36.689 ;
        RECT 28.186 36.671 36.558 36.735 ;
        RECT 28.14 36.717 36.512 36.781 ;
        RECT 28.094 36.763 36.466 36.827 ;
        RECT 28.048 36.809 36.42 36.873 ;
        RECT 28.002 36.855 36.374 36.919 ;
        RECT 27.956 36.901 36.328 36.965 ;
        RECT 27.91 36.947 36.282 37.011 ;
        RECT 27.864 36.993 36.236 37.057 ;
        RECT 27.818 37.039 36.19 37.103 ;
        RECT 27.772 37.085 36.144 37.149 ;
        RECT 27.726 37.131 36.098 37.195 ;
        RECT 27.68 37.177 36.052 37.241 ;
        RECT 27.634 37.223 36.006 37.287 ;
        RECT 27.588 37.269 35.96 37.333 ;
        RECT 27.542 37.315 35.914 37.379 ;
        RECT 27.496 37.361 35.868 37.425 ;
        RECT 27.45 37.407 35.822 37.471 ;
        RECT 27.404 37.453 35.776 37.517 ;
        RECT 27.358 37.499 35.73 37.563 ;
        RECT 27.312 37.545 35.684 37.609 ;
        RECT 27.266 37.591 35.638 37.655 ;
        RECT 27.22 37.637 35.592 37.701 ;
        RECT 27.174 37.683 35.546 37.747 ;
        RECT 27.128 37.729 35.5 37.793 ;
        RECT 27.082 37.775 35.454 37.839 ;
        RECT 27.036 37.821 35.408 37.885 ;
        RECT 26.99 37.867 35.362 37.931 ;
        RECT 26.944 37.913 35.316 37.977 ;
        RECT 26.898 37.959 35.27 38.023 ;
        RECT 26.852 38.005 35.224 38.069 ;
        RECT 26.806 38.051 35.178 38.115 ;
        RECT 26.76 38.097 35.132 38.161 ;
        RECT 26.714 38.143 35.086 38.207 ;
        RECT 26.668 38.189 35.04 38.253 ;
        RECT 26.622 38.235 34.994 38.299 ;
        RECT 26.576 38.281 34.948 38.345 ;
        RECT 26.53 38.327 34.902 38.391 ;
        RECT 26.484 38.373 34.856 38.437 ;
        RECT 26.438 38.419 34.81 38.483 ;
        RECT 26.392 38.465 34.764 38.529 ;
        RECT 26.346 38.511 34.718 38.575 ;
        RECT 26.3 38.557 34.672 38.621 ;
        RECT 26.254 38.603 34.626 38.667 ;
        RECT 26.208 38.649 34.58 38.713 ;
        RECT 26.162 38.695 34.534 38.759 ;
        RECT 26.116 38.741 34.488 38.805 ;
        RECT 26.07 38.787 34.442 38.851 ;
        RECT 26.024 38.833 34.396 38.897 ;
        RECT 25.978 38.879 34.35 38.943 ;
        RECT 25.932 38.925 34.304 38.989 ;
        RECT 25.886 38.971 34.258 39.035 ;
        RECT 25.84 39.017 34.212 39.081 ;
        RECT 25.794 39.063 34.166 39.127 ;
        RECT 25.748 39.109 34.12 39.173 ;
        RECT 25.702 39.155 34.074 39.219 ;
        RECT 25.656 39.201 34.028 39.265 ;
        RECT 25.61 39.247 33.982 39.311 ;
        RECT 25.564 39.293 33.936 39.357 ;
        RECT 25.518 39.339 33.89 39.403 ;
        RECT 25.472 39.385 33.844 39.449 ;
        RECT 25.426 39.431 33.798 39.495 ;
        RECT 25.38 39.477 33.752 39.541 ;
        RECT 25.334 39.523 33.706 39.587 ;
        RECT 25.288 39.569 33.66 39.633 ;
        RECT 25.242 39.615 33.614 39.679 ;
        RECT 25.196 39.661 33.568 39.725 ;
        RECT 25.15 39.707 33.522 39.771 ;
        RECT 25.104 39.753 33.476 39.817 ;
        RECT 25.058 39.799 33.43 39.863 ;
        RECT 25.012 39.845 33.384 39.909 ;
        RECT 24.966 39.891 33.338 39.955 ;
        RECT 24.92 39.937 33.292 40.001 ;
        RECT 24.874 39.983 33.246 40.047 ;
        RECT 24.828 40.029 33.2 40.093 ;
        RECT 24.782 40.075 33.154 40.139 ;
        RECT 24.736 40.121 33.108 40.185 ;
        RECT 24.69 40.167 33.062 40.231 ;
        RECT 24.644 40.213 33.016 40.277 ;
        RECT 24.598 40.259 32.97 40.323 ;
        RECT 24.552 40.305 32.924 40.369 ;
        RECT 24.506 40.351 32.878 40.415 ;
        RECT 24.46 40.397 32.832 40.461 ;
        RECT 24.414 40.443 32.786 40.507 ;
        RECT 24.368 40.489 32.74 40.553 ;
        RECT 24.322 40.535 32.694 40.599 ;
        RECT 24.276 40.581 32.648 40.645 ;
        RECT 24.23 40.627 32.602 40.691 ;
        RECT 24.184 40.673 32.556 40.737 ;
        RECT 24.138 40.719 32.51 40.783 ;
        RECT 24.092 40.765 32.464 40.829 ;
        RECT 24.046 40.811 32.418 40.875 ;
        RECT 24 40.857 32.372 40.921 ;
        RECT 23.954 40.903 32.326 40.967 ;
        RECT 23.908 40.949 32.28 41.013 ;
        RECT 23.862 40.995 32.234 41.059 ;
        RECT 23.816 41.041 32.188 41.105 ;
        RECT 23.77 41.087 32.142 41.151 ;
        RECT 23.724 41.133 32.096 41.197 ;
        RECT 23.678 41.179 32.05 41.243 ;
        RECT 23.632 41.225 32.004 41.289 ;
        RECT 23.586 41.271 31.958 41.335 ;
        RECT 23.54 41.317 31.912 41.381 ;
        RECT 23.494 41.363 31.866 41.427 ;
        RECT 23.448 41.409 31.82 41.473 ;
        RECT 23.402 41.455 31.774 41.519 ;
        RECT 23.356 41.501 31.728 41.565 ;
        RECT 23.31 41.547 31.682 41.611 ;
        RECT 23.264 41.593 31.636 41.657 ;
        RECT 23.218 41.639 31.59 41.703 ;
        RECT 23.172 41.685 31.544 41.749 ;
        RECT 23.126 41.731 31.498 41.795 ;
        RECT 23.08 41.777 31.452 41.841 ;
        RECT 23.034 41.823 31.406 41.887 ;
        RECT 22.988 41.869 31.36 41.933 ;
        RECT 22.942 41.915 31.314 41.979 ;
        RECT 22.896 41.961 31.268 42.025 ;
        RECT 22.85 42.007 31.222 42.071 ;
        RECT 22.804 42.053 31.176 42.117 ;
        RECT 22.758 42.099 31.13 42.163 ;
        RECT 22.712 42.145 31.084 42.209 ;
        RECT 22.666 42.191 31.038 42.255 ;
        RECT 22.62 42.237 30.992 42.301 ;
        RECT 22.574 42.283 30.946 42.347 ;
        RECT 22.528 42.329 30.9 42.393 ;
        RECT 22.482 42.375 30.854 42.439 ;
        RECT 22.436 42.421 30.808 42.485 ;
        RECT 22.39 42.467 30.762 42.531 ;
        RECT 22.344 42.513 30.716 42.577 ;
        RECT 22.298 42.559 30.67 42.623 ;
        RECT 22.252 42.605 30.624 42.669 ;
        RECT 22.206 42.651 30.578 42.715 ;
        RECT 22.16 42.697 30.532 42.761 ;
        RECT 22.114 42.743 30.486 42.807 ;
        RECT 22.068 42.789 30.44 42.853 ;
        RECT 22.022 42.835 30.394 42.899 ;
        RECT 21.976 42.881 30.348 42.945 ;
        RECT 21.93 42.927 30.302 42.991 ;
        RECT 21.884 42.973 30.256 43.037 ;
        RECT 21.838 43.019 30.21 43.083 ;
        RECT 21.792 43.065 30.164 43.129 ;
        RECT 21.746 43.111 30.118 43.175 ;
        RECT 21.7 43.157 30.072 43.221 ;
        RECT 21.654 43.203 30.026 43.267 ;
        RECT 21.608 43.249 29.98 43.313 ;
        RECT 21.562 43.295 29.934 43.359 ;
        RECT 21.516 43.341 29.888 43.405 ;
        RECT 21.47 43.387 29.842 43.451 ;
        RECT 21.424 43.433 29.796 43.497 ;
        RECT 21.378 43.479 29.75 43.543 ;
        RECT 21.332 43.525 29.704 43.589 ;
        RECT 21.286 43.571 29.658 43.635 ;
        RECT 21.24 43.617 29.612 43.681 ;
        RECT 21.194 43.663 29.566 43.727 ;
        RECT 21.148 43.709 29.52 43.773 ;
        RECT 21.102 43.755 29.474 43.819 ;
        RECT 21.056 43.801 29.428 43.865 ;
        RECT 21.01 43.847 29.382 43.911 ;
        RECT 20.964 43.893 29.336 43.957 ;
        RECT 20.918 43.939 29.29 44.003 ;
        RECT 20.872 43.985 29.244 44.049 ;
        RECT 20.826 44.031 29.198 44.095 ;
        RECT 20.78 44.077 29.152 44.141 ;
        RECT 20.734 44.123 29.106 44.187 ;
        RECT 20.688 44.169 29.06 44.233 ;
        RECT 20.642 44.215 29.014 44.279 ;
        RECT 20.596 44.261 28.968 44.325 ;
        RECT 20.55 44.307 28.922 44.371 ;
        RECT 20.504 44.353 28.876 44.417 ;
        RECT 20.458 44.399 28.83 44.463 ;
        RECT 20.412 44.445 28.784 44.509 ;
        RECT 20.366 44.491 28.738 44.555 ;
        RECT 20.32 44.537 28.692 44.601 ;
        RECT 20.274 44.583 28.646 44.647 ;
        RECT 20.228 44.629 28.6 44.693 ;
        RECT 20.182 44.675 28.554 44.739 ;
        RECT 20.136 44.721 28.508 44.785 ;
        RECT 20.09 44.767 28.462 44.831 ;
        RECT 20.044 44.813 28.416 44.877 ;
        RECT 19.998 44.859 28.37 44.923 ;
        RECT 19.952 44.905 28.324 44.969 ;
        RECT 19.906 44.951 28.278 45.015 ;
        RECT 19.86 44.997 28.232 45.061 ;
        RECT 19.814 45.043 28.186 45.107 ;
        RECT 19.768 45.089 28.14 45.153 ;
        RECT 19.722 45.135 28.094 45.199 ;
        RECT 19.676 45.181 28.048 45.245 ;
        RECT 19.63 45.227 28.002 45.291 ;
        RECT 19.584 45.273 27.956 45.337 ;
        RECT 19.538 45.319 27.91 45.383 ;
        RECT 19.492 45.365 27.864 45.429 ;
        RECT 19.446 45.411 27.818 45.475 ;
        RECT 19.4 45.457 27.772 45.521 ;
        RECT 19.354 45.503 27.726 45.567 ;
        RECT 19.308 45.549 27.68 45.613 ;
        RECT 19.262 45.595 27.634 45.659 ;
        RECT 19.216 45.641 27.588 45.705 ;
        RECT 19.17 45.687 27.542 45.751 ;
        RECT 19.124 45.733 27.496 45.797 ;
        RECT 19.078 45.779 27.45 45.843 ;
        RECT 19.032 45.825 27.404 45.889 ;
        RECT 18.986 45.871 27.358 45.935 ;
        RECT 18.94 45.917 27.312 45.981 ;
        RECT 18.894 45.963 27.266 46.027 ;
        RECT 18.848 46.009 27.22 46.073 ;
        RECT 18.802 46.055 27.174 46.119 ;
        RECT 18.756 46.101 27.128 46.165 ;
        RECT 18.71 46.147 27.082 46.211 ;
        RECT 18.664 46.193 27.036 46.257 ;
        RECT 18.618 46.239 26.99 46.303 ;
        RECT 18.572 46.285 26.944 46.349 ;
        RECT 18.526 46.331 26.898 46.395 ;
        RECT 18.48 46.377 26.852 46.441 ;
        RECT 18.434 46.423 26.806 46.487 ;
        RECT 18.388 46.469 26.76 46.533 ;
        RECT 18.342 46.515 26.714 46.579 ;
        RECT 18.296 46.561 26.668 46.625 ;
        RECT 18.25 46.607 26.622 46.671 ;
        RECT 18.204 46.653 26.576 46.717 ;
        RECT 18.158 46.699 26.53 46.763 ;
        RECT 18.112 46.745 26.484 46.809 ;
        RECT 18.066 46.791 26.438 46.855 ;
        RECT 18.02 46.837 26.392 46.901 ;
        RECT 17.974 46.883 26.346 46.947 ;
        RECT 17.928 46.929 26.3 46.993 ;
        RECT 17.882 46.975 26.254 47.039 ;
        RECT 17.836 47.021 26.208 47.085 ;
        RECT 17.79 47.067 26.162 47.131 ;
        RECT 17.744 47.113 26.116 47.177 ;
        RECT 17.698 47.159 26.07 47.223 ;
        RECT 17.652 47.205 26.024 47.269 ;
        RECT 17.606 47.251 25.978 47.315 ;
        RECT 17.56 47.297 25.932 47.361 ;
        RECT 17.514 47.343 25.886 47.407 ;
        RECT 17.468 47.389 25.84 47.453 ;
        RECT 17.422 47.435 25.794 47.499 ;
        RECT 17.376 47.481 25.748 47.545 ;
        RECT 17.33 47.527 25.702 47.591 ;
        RECT 17.284 47.573 25.656 47.637 ;
        RECT 17.238 47.619 25.61 47.683 ;
        RECT 17.192 47.665 25.564 47.729 ;
        RECT 17.146 47.711 25.518 47.775 ;
        RECT 17.1 47.757 25.472 47.821 ;
        RECT 17.054 47.803 25.426 47.867 ;
        RECT 17.008 47.849 25.38 47.913 ;
        RECT 16.962 47.895 25.334 47.959 ;
        RECT 16.916 47.941 25.288 48.005 ;
        RECT 16.87 47.987 25.242 48.051 ;
        RECT 16.824 48.033 25.196 48.097 ;
        RECT 16.778 48.079 25.15 48.143 ;
        RECT 16.732 48.125 25.104 48.189 ;
        RECT 16.686 48.171 25.058 48.235 ;
        RECT 16.64 48.217 25.012 48.281 ;
        RECT 16.594 48.263 24.966 48.327 ;
        RECT 16.548 48.309 24.92 48.373 ;
        RECT 16.502 48.355 24.874 48.419 ;
        RECT 16.456 48.401 24.828 48.465 ;
        RECT 16.41 48.447 24.782 48.511 ;
        RECT 16.364 48.493 24.736 48.557 ;
        RECT 16.318 48.539 24.69 48.603 ;
        RECT 16.272 48.585 24.644 48.649 ;
        RECT 16.226 48.631 24.598 48.695 ;
        RECT 16.18 48.677 24.552 48.741 ;
        RECT 16.134 48.723 24.506 48.787 ;
        RECT 16.088 48.769 24.46 48.833 ;
        RECT 16.042 48.815 24.414 48.879 ;
        RECT 15.996 48.861 24.368 48.925 ;
        RECT 15.95 48.907 24.322 48.971 ;
        RECT 15.904 48.953 24.276 49.017 ;
        RECT 15.858 48.999 24.23 49.063 ;
        RECT 15.812 49.045 24.184 49.109 ;
        RECT 15.766 49.091 24.138 49.155 ;
        RECT 15.72 49.137 24.092 49.201 ;
        RECT 15.674 49.183 24.046 49.247 ;
        RECT 15.628 49.229 24 49.293 ;
        RECT 15.582 49.275 23.954 49.339 ;
        RECT 15.536 49.321 23.908 49.385 ;
        RECT 15.49 49.367 23.862 49.431 ;
        RECT 15.444 49.413 23.816 49.477 ;
        RECT 15.398 49.459 23.77 49.523 ;
        RECT 15.352 49.505 23.724 49.569 ;
        RECT 15.306 49.551 23.678 49.615 ;
        RECT 15.26 49.597 23.632 49.661 ;
        RECT 15.214 49.643 23.586 49.707 ;
        RECT 15.168 49.689 23.54 49.753 ;
        RECT 15.122 49.735 23.494 49.799 ;
        RECT 15.076 49.781 23.448 49.845 ;
        RECT 15.03 49.827 23.402 49.891 ;
        RECT 14.984 49.873 23.356 49.937 ;
        RECT 14.938 49.919 23.31 49.983 ;
        RECT 14.892 49.965 23.264 50.029 ;
        RECT 14.846 50.011 23.218 50.075 ;
        RECT 14.8 50.057 23.172 50.121 ;
        RECT 14.754 50.103 23.126 50.167 ;
        RECT 14.708 50.149 23.08 50.213 ;
        RECT 14.662 50.195 23.034 50.259 ;
        RECT 14.616 50.241 22.988 50.305 ;
        RECT 14.57 50.287 22.942 50.351 ;
        RECT 14.524 50.333 22.896 50.397 ;
        RECT 14.478 50.379 22.85 50.443 ;
        RECT 14.432 50.425 22.804 50.489 ;
        RECT 14.386 50.471 22.758 50.535 ;
        RECT 14.34 50.517 22.712 50.581 ;
        RECT 14.294 50.563 22.666 50.627 ;
        RECT 14.248 50.609 22.62 50.673 ;
        RECT 14.202 50.655 22.574 50.719 ;
        RECT 14.156 50.701 22.528 50.765 ;
        RECT 14.11 50.747 22.482 50.811 ;
        RECT 14.064 50.793 22.436 50.857 ;
        RECT 14.018 50.839 22.39 50.903 ;
        RECT 13.972 50.885 22.344 50.949 ;
        RECT 13.926 50.931 22.298 50.995 ;
        RECT 13.88 50.977 22.252 51.041 ;
        RECT 13.834 51.023 22.206 51.087 ;
        RECT 13.788 51.069 22.16 51.133 ;
        RECT 13.742 51.115 22.114 51.179 ;
        RECT 13.696 51.161 22.068 51.225 ;
        RECT 13.65 51.207 22.022 51.271 ;
        RECT 13.604 51.253 21.976 51.317 ;
        RECT 13.558 51.299 21.93 51.363 ;
    END
    PORT
      LAYER QB ;
        RECT 67.73 42.6 80 47.4 ;
        RECT 62.902 47.405 69.708 47.435 ;
        RECT 60.97 49.337 67.73 49.412 ;
        RECT 61.016 49.291 67.776 49.367 ;
        RECT 67.686 42.622 67.73 49.412 ;
        RECT 60.924 49.383 67.686 49.457 ;
        RECT 61.062 49.245 67.822 49.321 ;
        RECT 67.64 42.667 67.686 49.457 ;
        RECT 60.878 49.429 67.64 49.503 ;
        RECT 61.108 49.199 67.868 49.275 ;
        RECT 67.594 42.713 67.64 49.503 ;
        RECT 60.832 49.475 67.594 49.549 ;
        RECT 61.154 49.153 67.914 49.229 ;
        RECT 67.548 42.759 67.594 49.549 ;
        RECT 60.786 49.521 67.548 49.595 ;
        RECT 61.2 49.107 67.96 49.183 ;
        RECT 67.502 42.805 67.548 49.595 ;
        RECT 60.74 49.567 67.502 49.641 ;
        RECT 61.246 49.061 68.006 49.137 ;
        RECT 67.456 42.851 67.502 49.641 ;
        RECT 60.694 49.613 67.456 49.687 ;
        RECT 61.292 49.015 68.052 49.091 ;
        RECT 67.41 42.897 67.456 49.687 ;
        RECT 60.648 49.659 67.41 49.733 ;
        RECT 61.338 48.969 68.098 49.045 ;
        RECT 67.364 42.943 67.41 49.733 ;
        RECT 60.602 49.705 67.364 49.779 ;
        RECT 61.384 48.923 68.144 48.999 ;
        RECT 67.318 42.989 67.364 49.779 ;
        RECT 60.556 49.751 67.318 49.825 ;
        RECT 61.43 48.877 68.19 48.953 ;
        RECT 67.272 43.035 67.318 49.825 ;
        RECT 60.51 49.797 67.272 49.871 ;
        RECT 61.476 48.831 68.236 48.907 ;
        RECT 67.226 43.081 67.272 49.871 ;
        RECT 60.464 49.843 67.226 49.917 ;
        RECT 61.522 48.785 68.282 48.861 ;
        RECT 67.18 43.127 67.226 49.917 ;
        RECT 60.418 49.889 67.18 49.963 ;
        RECT 61.568 48.739 68.328 48.815 ;
        RECT 67.134 43.173 67.18 49.963 ;
        RECT 60.372 49.935 67.134 50.009 ;
        RECT 61.614 48.693 68.374 48.769 ;
        RECT 67.088 43.219 67.134 50.009 ;
        RECT 60.326 49.981 67.088 50.055 ;
        RECT 61.66 48.647 68.42 48.723 ;
        RECT 67.042 43.265 67.088 50.055 ;
        RECT 60.28 50.027 67.042 50.101 ;
        RECT 61.706 48.601 68.466 48.677 ;
        RECT 66.996 43.311 67.042 50.101 ;
        RECT 60.234 50.073 66.996 50.147 ;
        RECT 61.752 48.555 68.512 48.631 ;
        RECT 66.95 43.357 66.996 50.147 ;
        RECT 60.188 50.119 66.95 50.193 ;
        RECT 61.798 48.509 68.558 48.585 ;
        RECT 66.904 43.403 66.95 50.193 ;
        RECT 60.142 50.165 66.904 50.239 ;
        RECT 61.844 48.463 68.604 48.539 ;
        RECT 66.858 43.449 66.904 50.239 ;
        RECT 60.096 50.211 66.858 50.285 ;
        RECT 61.89 48.417 68.65 48.493 ;
        RECT 66.812 43.495 66.858 50.285 ;
        RECT 60.05 50.257 66.812 50.331 ;
        RECT 61.936 48.371 68.696 48.447 ;
        RECT 66.766 43.541 66.812 50.331 ;
        RECT 60.004 50.303 66.766 50.377 ;
        RECT 61.982 48.325 68.742 48.401 ;
        RECT 66.72 43.587 66.766 50.377 ;
        RECT 59.958 50.349 66.72 50.423 ;
        RECT 62.028 48.279 68.788 48.355 ;
        RECT 66.674 43.633 66.72 50.423 ;
        RECT 59.912 50.395 66.674 50.469 ;
        RECT 62.074 48.233 68.834 48.309 ;
        RECT 66.628 43.679 66.674 50.469 ;
        RECT 59.866 50.441 66.628 50.515 ;
        RECT 62.12 48.187 68.88 48.263 ;
        RECT 66.582 43.725 66.628 50.515 ;
        RECT 59.82 50.487 66.582 50.561 ;
        RECT 62.166 48.141 68.926 48.217 ;
        RECT 66.536 43.771 66.582 50.561 ;
        RECT 59.774 50.533 66.536 50.607 ;
        RECT 62.212 48.095 68.972 48.171 ;
        RECT 66.49 43.817 66.536 50.607 ;
        RECT 59.728 50.579 66.49 50.653 ;
        RECT 62.258 48.049 69.018 48.125 ;
        RECT 66.444 43.863 66.49 50.653 ;
        RECT 59.682 50.625 66.444 50.699 ;
        RECT 62.304 48.003 69.064 48.079 ;
        RECT 66.398 43.909 66.444 50.699 ;
        RECT 59.636 50.671 66.398 50.745 ;
        RECT 62.35 47.957 69.11 48.033 ;
        RECT 66.352 43.955 66.398 50.745 ;
        RECT 59.59 50.717 66.352 50.791 ;
        RECT 62.396 47.911 69.156 47.987 ;
        RECT 66.306 44.001 66.352 50.791 ;
        RECT 59.544 50.763 66.306 50.837 ;
        RECT 62.442 47.865 69.202 47.941 ;
        RECT 66.26 44.047 66.306 50.837 ;
        RECT 59.498 50.809 66.26 50.883 ;
        RECT 62.488 47.819 69.248 47.895 ;
        RECT 66.214 44.093 66.26 50.883 ;
        RECT 59.452 50.855 66.214 50.929 ;
        RECT 62.534 47.773 69.294 47.849 ;
        RECT 66.168 44.139 66.214 50.929 ;
        RECT 59.406 50.901 66.168 50.975 ;
        RECT 62.58 47.727 69.34 47.803 ;
        RECT 66.122 44.185 66.168 50.975 ;
        RECT 59.36 50.947 66.122 51.021 ;
        RECT 62.626 47.681 69.386 47.757 ;
        RECT 66.076 44.231 66.122 51.021 ;
        RECT 59.314 50.993 66.076 51.067 ;
        RECT 62.672 47.635 69.432 47.711 ;
        RECT 66.03 44.277 66.076 51.067 ;
        RECT 59.268 51.039 66.03 51.113 ;
        RECT 62.718 47.589 69.478 47.665 ;
        RECT 65.984 44.323 66.03 51.113 ;
        RECT 59.222 51.085 65.984 51.159 ;
        RECT 62.764 47.543 69.524 47.619 ;
        RECT 65.938 44.369 65.984 51.159 ;
        RECT 59.176 51.131 65.938 51.205 ;
        RECT 62.81 47.497 69.57 47.573 ;
        RECT 65.892 44.415 65.938 51.205 ;
        RECT 59.13 51.177 65.892 51.251 ;
        RECT 62.856 47.451 69.616 47.527 ;
        RECT 65.846 44.461 65.892 51.251 ;
        RECT 59.084 51.223 65.846 51.297 ;
        RECT 62.902 47.405 69.662 47.481 ;
        RECT 65.8 44.507 65.846 51.297 ;
        RECT 59.038 51.269 65.8 51.343 ;
        RECT 62.948 47.359 69.72 47.406 ;
        RECT 65.754 44.553 65.8 51.343 ;
        RECT 58.992 51.315 65.754 51.389 ;
        RECT 62.994 47.313 80 47.4 ;
        RECT 65.708 44.599 65.754 51.389 ;
        RECT 58.946 51.361 65.708 51.435 ;
        RECT 63.04 47.267 80 47.4 ;
        RECT 65.662 44.645 65.708 51.435 ;
        RECT 58.9 51.407 65.662 51.481 ;
        RECT 63.086 47.221 80 47.4 ;
        RECT 65.616 44.691 65.662 51.481 ;
        RECT 58.854 51.453 65.616 51.527 ;
        RECT 63.132 47.175 80 47.4 ;
        RECT 65.57 44.737 65.616 51.527 ;
        RECT 58.808 51.499 65.57 51.573 ;
        RECT 63.178 47.129 80 47.4 ;
        RECT 65.524 44.783 65.57 51.573 ;
        RECT 58.762 51.545 65.524 51.619 ;
        RECT 63.224 47.083 80 47.4 ;
        RECT 65.478 44.829 65.524 51.619 ;
        RECT 58.716 51.591 65.478 51.665 ;
        RECT 63.27 47.037 80 47.4 ;
        RECT 65.432 44.875 65.478 51.665 ;
        RECT 58.67 51.637 65.432 51.711 ;
        RECT 63.316 46.991 80 47.4 ;
        RECT 65.386 44.921 65.432 51.711 ;
        RECT 58.624 51.683 65.386 51.757 ;
        RECT 63.362 46.945 80 47.4 ;
        RECT 65.34 44.967 65.386 51.757 ;
        RECT 58.578 51.729 65.34 51.803 ;
        RECT 63.408 46.899 80 47.4 ;
        RECT 65.294 45.013 65.34 51.803 ;
        RECT 58.532 51.775 65.294 51.849 ;
        RECT 63.454 46.853 80 47.4 ;
        RECT 65.248 45.059 65.294 51.849 ;
        RECT 58.486 51.821 65.248 51.895 ;
        RECT 63.5 46.807 80 47.4 ;
        RECT 65.202 45.105 65.248 51.895 ;
        RECT 58.44 51.867 65.202 51.941 ;
        RECT 63.546 46.761 80 47.4 ;
        RECT 65.156 45.151 65.202 51.941 ;
        RECT 58.394 51.913 65.156 51.987 ;
        RECT 63.592 46.715 80 47.4 ;
        RECT 65.11 45.197 65.156 51.987 ;
        RECT 58.348 51.959 65.11 52.033 ;
        RECT 63.638 46.669 80 47.4 ;
        RECT 65.064 45.243 65.11 52.033 ;
        RECT 58.302 52.005 65.064 52.079 ;
        RECT 63.684 46.623 80 47.4 ;
        RECT 65.018 45.289 65.064 52.079 ;
        RECT 58.256 52.051 65.018 52.125 ;
        RECT 63.73 46.577 80 47.4 ;
        RECT 64.972 45.335 65.018 52.125 ;
        RECT 58.21 52.097 64.972 52.171 ;
        RECT 63.776 46.531 80 47.4 ;
        RECT 64.926 45.381 64.972 52.171 ;
        RECT 58.164 52.143 64.926 52.217 ;
        RECT 63.822 46.485 80 47.4 ;
        RECT 64.88 45.427 64.926 52.217 ;
        RECT 58.118 52.189 64.88 52.263 ;
        RECT 63.868 46.439 80 47.4 ;
        RECT 64.834 45.473 64.88 52.263 ;
        RECT 58.072 52.235 64.834 52.309 ;
        RECT 63.914 46.393 80 47.4 ;
        RECT 64.788 45.519 64.834 52.309 ;
        RECT 58.026 52.281 64.788 52.355 ;
        RECT 63.96 46.347 80 47.4 ;
        RECT 64.742 45.565 64.788 52.355 ;
        RECT 57.98 52.327 64.742 52.401 ;
        RECT 64.006 46.301 80 47.4 ;
        RECT 64.696 45.611 64.742 52.401 ;
        RECT 57.934 52.373 64.696 52.447 ;
        RECT 64.052 46.255 80 47.4 ;
        RECT 64.65 45.657 64.696 52.447 ;
        RECT 57.888 52.419 64.65 52.493 ;
        RECT 64.098 46.209 80 47.4 ;
        RECT 64.604 45.703 64.65 52.493 ;
        RECT 57.842 52.465 64.604 52.539 ;
        RECT 64.144 46.163 80 47.4 ;
        RECT 64.558 45.749 64.604 52.539 ;
        RECT 57.796 52.511 64.558 52.585 ;
        RECT 64.19 46.117 80 47.4 ;
        RECT 64.512 45.795 64.558 52.585 ;
        RECT 57.75 52.557 64.512 52.631 ;
        RECT 64.236 46.071 80 47.4 ;
        RECT 64.466 45.841 64.512 52.631 ;
        RECT 57.704 52.603 64.466 52.677 ;
        RECT 64.282 46.025 80 47.4 ;
        RECT 64.42 45.887 64.466 52.677 ;
        RECT 57.658 52.649 64.42 52.723 ;
        RECT 64.328 45.979 80 47.4 ;
        RECT 64.374 45.933 64.42 52.723 ;
        RECT 57.612 52.695 64.374 52.769 ;
        RECT 57.566 52.741 64.328 52.815 ;
        RECT 57.52 52.787 64.282 52.861 ;
        RECT 57.474 52.833 64.236 52.907 ;
        RECT 57.428 52.879 64.19 52.953 ;
        RECT 57.382 52.925 64.144 52.999 ;
        RECT 57.336 52.971 64.098 53.045 ;
        RECT 57.29 53.017 64.052 53.091 ;
        RECT 57.244 53.063 64.006 53.137 ;
        RECT 57.198 53.109 63.96 53.183 ;
        RECT 57.152 53.155 63.914 53.229 ;
        RECT 57.106 53.201 63.868 53.275 ;
        RECT 57.06 53.247 63.822 53.321 ;
        RECT 57.014 53.293 63.776 53.367 ;
        RECT 56.968 53.339 63.73 53.413 ;
        RECT 56.922 53.385 63.684 53.459 ;
        RECT 56.876 53.431 63.638 53.505 ;
        RECT 56.83 53.477 63.592 53.551 ;
        RECT 56.784 53.523 63.546 53.597 ;
        RECT 56.738 53.569 63.5 53.643 ;
        RECT 56.692 53.615 63.454 53.689 ;
        RECT 56.646 53.661 63.408 53.735 ;
        RECT 56.6 53.707 63.362 53.781 ;
        RECT 56.554 53.753 63.316 53.827 ;
        RECT 56.508 53.799 63.27 53.873 ;
        RECT 56.462 53.845 63.224 53.919 ;
        RECT 56.416 53.891 63.178 53.965 ;
        RECT 56.37 53.937 63.132 54.011 ;
        RECT 56.324 53.983 63.086 54.057 ;
        RECT 56.278 54.029 63.04 54.103 ;
        RECT 56.232 54.075 62.994 54.149 ;
        RECT 56.186 54.121 62.948 54.195 ;
        RECT 56.14 54.167 62.902 54.241 ;
        RECT 56.094 54.213 62.856 54.287 ;
        RECT 56.048 54.259 62.81 54.333 ;
        RECT 56.002 54.305 62.764 54.379 ;
        RECT 55.956 54.351 62.718 54.425 ;
        RECT 55.91 54.397 62.672 54.471 ;
        RECT 55.864 54.443 62.626 54.517 ;
        RECT 55.818 54.489 62.58 54.563 ;
        RECT 55.772 54.535 62.534 54.609 ;
        RECT 55.726 54.581 62.488 54.655 ;
        RECT 55.68 54.627 62.442 54.701 ;
        RECT 55.634 54.673 62.396 54.747 ;
        RECT 55.588 54.719 62.35 54.793 ;
        RECT 55.542 54.765 62.304 54.839 ;
        RECT 55.496 54.811 62.258 54.885 ;
        RECT 55.45 54.857 62.212 54.931 ;
        RECT 55.404 54.903 62.166 54.977 ;
        RECT 55.358 54.949 62.12 55.023 ;
        RECT 55.312 54.995 62.074 55.069 ;
        RECT 55.266 55.041 62.028 55.115 ;
        RECT 55.22 55.087 61.982 55.161 ;
        RECT 55.174 55.133 61.936 55.207 ;
        RECT 55.128 55.179 61.89 55.253 ;
        RECT 55.082 55.225 61.844 55.299 ;
        RECT 55.036 55.271 61.798 55.345 ;
        RECT 54.99 55.317 61.752 55.391 ;
        RECT 54.944 55.363 61.706 55.437 ;
        RECT 54.898 55.409 61.66 55.483 ;
        RECT 54.852 55.455 61.614 55.529 ;
        RECT 54.806 55.501 61.568 55.575 ;
        RECT 54.76 55.547 61.522 55.621 ;
        RECT 54.714 55.593 61.476 55.667 ;
        RECT 54.668 55.639 61.43 55.713 ;
        RECT 54.622 55.685 61.384 55.759 ;
        RECT 54.576 55.731 61.338 55.805 ;
        RECT 54.53 55.777 61.292 55.851 ;
        RECT 54.484 55.823 61.246 55.897 ;
        RECT 54.438 55.869 61.2 55.943 ;
        RECT 54.392 55.915 61.154 55.989 ;
        RECT 54.346 55.961 61.108 56.035 ;
        RECT 54.3 56.007 61.062 56.081 ;
        RECT 54.254 56.053 61.016 56.127 ;
        RECT 54.208 56.099 60.97 56.173 ;
        RECT 54.162 56.145 60.924 56.219 ;
        RECT 54.116 56.191 60.878 56.265 ;
        RECT 54.07 56.237 60.832 56.311 ;
        RECT 54.024 56.283 60.786 56.357 ;
        RECT 53.978 56.329 60.74 56.403 ;
        RECT 53.932 56.375 60.694 56.449 ;
        RECT 53.886 56.421 60.648 56.495 ;
        RECT 53.84 56.467 60.602 56.541 ;
        RECT 53.794 56.513 60.556 56.587 ;
        RECT 53.748 56.559 60.51 56.633 ;
        RECT 53.702 56.605 60.464 56.679 ;
        RECT 53.656 56.651 60.418 56.725 ;
        RECT 53.61 56.697 60.372 56.771 ;
        RECT 53.564 56.743 60.326 56.817 ;
        RECT 53.518 56.789 60.28 56.863 ;
        RECT 53.472 56.835 60.234 56.909 ;
        RECT 53.426 56.881 60.188 56.955 ;
        RECT 53.38 56.927 60.142 57.001 ;
        RECT 53.334 56.973 60.096 57.047 ;
        RECT 53.288 57.019 60.05 57.093 ;
        RECT 53.242 57.065 60.004 57.139 ;
        RECT 53.196 57.111 59.958 57.185 ;
        RECT 53.15 57.157 59.912 57.231 ;
        RECT 53.104 57.203 59.866 57.277 ;
        RECT 53.058 57.249 59.82 57.323 ;
        RECT 53.012 57.295 59.774 57.369 ;
        RECT 52.966 57.341 59.728 57.415 ;
        RECT 52.92 57.387 59.682 57.461 ;
        RECT 52.874 57.433 59.636 57.507 ;
        RECT 52.828 57.479 59.59 57.553 ;
        RECT 52.782 57.525 59.544 57.599 ;
        RECT 52.736 57.571 59.498 57.645 ;
        RECT 52.69 57.617 59.452 57.691 ;
        RECT 52.644 57.663 59.406 57.737 ;
        RECT 52.598 57.709 59.36 57.783 ;
        RECT 52.552 57.755 59.314 57.829 ;
        RECT 52.506 57.801 59.268 57.875 ;
        RECT 52.46 57.847 59.222 57.921 ;
        RECT 52.414 57.893 59.176 57.967 ;
        RECT 52.368 57.939 59.13 58.013 ;
        RECT 52.322 57.985 59.084 58.059 ;
        RECT 52.276 58.031 59.038 58.105 ;
        RECT 52.23 58.077 58.992 58.151 ;
        RECT 52.184 58.123 58.946 58.197 ;
        RECT 52.138 58.169 58.9 58.243 ;
        RECT 52.092 58.215 58.854 58.289 ;
        RECT 52.046 58.261 58.808 58.335 ;
        RECT 52 58.307 58.762 58.381 ;
        RECT 51.954 58.353 58.716 58.427 ;
        RECT 51.908 58.399 58.67 58.473 ;
        RECT 51.862 58.445 58.624 58.519 ;
        RECT 51.816 58.491 58.578 58.565 ;
        RECT 51.77 58.537 58.532 58.611 ;
        RECT 51.724 58.583 58.486 58.657 ;
        RECT 51.678 58.629 58.44 58.703 ;
        RECT 51.632 58.675 58.394 58.749 ;
        RECT 51.586 58.721 58.348 58.795 ;
        RECT 51.54 58.767 58.302 58.841 ;
        RECT 51.494 58.813 58.256 58.887 ;
        RECT 51.448 58.859 58.21 58.933 ;
        RECT 51.402 58.905 58.164 58.979 ;
        RECT 51.356 58.951 58.118 59.025 ;
        RECT 51.31 58.997 58.072 59.071 ;
        RECT 51.264 59.043 58.026 59.117 ;
        RECT 51.218 59.089 57.98 59.163 ;
        RECT 51.172 59.135 57.934 59.209 ;
        RECT 51.126 59.181 57.888 59.255 ;
        RECT 51.08 59.227 57.842 59.301 ;
        RECT 51.034 59.273 57.796 59.347 ;
        RECT 50.988 59.319 57.75 59.393 ;
        RECT 50.942 59.365 57.704 59.439 ;
        RECT 50.896 59.411 57.658 59.485 ;
        RECT 50.85 59.457 57.612 59.531 ;
        RECT 50.804 59.503 57.566 59.577 ;
        RECT 50.758 59.549 57.52 59.623 ;
        RECT 50.712 59.595 57.474 59.669 ;
        RECT 50.666 59.641 57.428 59.715 ;
        RECT 50.62 59.687 57.382 59.761 ;
        RECT 50.574 59.733 57.336 59.807 ;
        RECT 50.528 59.779 57.29 59.853 ;
        RECT 50.482 59.825 57.244 59.899 ;
        RECT 50.436 59.871 57.198 59.945 ;
        RECT 50.39 59.917 57.152 59.991 ;
        RECT 50.344 59.963 57.106 60.037 ;
        RECT 50.298 60.009 57.06 60.083 ;
        RECT 50.252 60.055 57.014 60.129 ;
        RECT 50.206 60.101 56.968 60.175 ;
        RECT 50.16 60.147 56.922 60.221 ;
        RECT 50.114 60.193 56.876 60.267 ;
        RECT 50.068 60.239 56.83 60.313 ;
        RECT 50.022 60.285 56.784 60.359 ;
        RECT 49.976 60.331 56.738 60.405 ;
        RECT 49.93 60.377 56.692 60.451 ;
        RECT 49.884 60.423 56.646 60.497 ;
        RECT 49.838 60.469 56.6 60.543 ;
        RECT 49.792 60.515 56.554 60.589 ;
        RECT 49.746 60.561 56.508 60.635 ;
        RECT 49.7 60.607 56.462 60.681 ;
        RECT 49.654 60.653 56.416 60.727 ;
        RECT 49.608 60.699 56.37 60.773 ;
        RECT 49.562 60.745 56.324 60.819 ;
        RECT 49.516 60.791 56.278 60.865 ;
        RECT 49.47 60.837 56.232 60.911 ;
        RECT 49.424 60.883 56.186 60.957 ;
        RECT 49.378 60.929 56.14 61.003 ;
        RECT 49.332 60.975 56.094 61.049 ;
        RECT 49.286 61.021 56.048 61.095 ;
        RECT 49.24 61.067 56.002 61.141 ;
        RECT 49.194 61.113 55.956 61.187 ;
        RECT 49.148 61.159 55.91 61.233 ;
        RECT 49.102 61.205 55.864 61.279 ;
        RECT 49.056 61.251 55.818 61.325 ;
        RECT 49.01 61.297 55.772 61.371 ;
        RECT 48.964 61.343 55.726 61.417 ;
        RECT 48.918 61.389 55.68 61.463 ;
        RECT 48.872 61.435 55.634 61.509 ;
        RECT 48.826 61.481 55.588 61.555 ;
        RECT 48.78 61.527 55.542 61.601 ;
        RECT 48.734 61.573 55.496 61.647 ;
        RECT 48.688 61.619 55.45 61.693 ;
        RECT 48.642 61.665 55.404 61.739 ;
        RECT 48.596 61.711 55.358 61.785 ;
        RECT 48.55 61.757 55.312 61.831 ;
        RECT 48.504 61.803 55.266 61.877 ;
        RECT 48.458 61.849 55.22 61.923 ;
        RECT 48.412 61.895 55.174 61.969 ;
        RECT 48.366 61.941 55.128 62.015 ;
        RECT 48.32 61.987 55.082 62.061 ;
        RECT 48.274 62.033 55.036 62.107 ;
        RECT 48.228 62.079 54.99 62.153 ;
        RECT 48.182 62.125 54.944 62.199 ;
        RECT 48.136 62.171 54.898 62.245 ;
        RECT 48.09 62.217 54.852 62.291 ;
        RECT 48.044 62.263 54.806 62.337 ;
        RECT 47.998 62.309 54.76 62.383 ;
        RECT 47.952 62.355 54.714 62.429 ;
        RECT 47.906 62.401 54.668 62.475 ;
        RECT 47.86 62.447 54.622 62.521 ;
        RECT 47.814 62.493 54.576 62.567 ;
        RECT 47.768 62.539 54.53 62.613 ;
        RECT 47.722 62.585 54.484 62.659 ;
        RECT 47.676 62.631 54.438 62.705 ;
        RECT 47.63 62.677 54.392 62.751 ;
        RECT 47.584 62.723 54.346 62.797 ;
        RECT 47.538 62.769 54.3 62.843 ;
        RECT 47.492 62.815 54.254 62.889 ;
        RECT 47.446 62.861 54.208 62.935 ;
        RECT 47.384 62.938 54.162 62.981 ;
        RECT 47.4 62.907 54.162 62.981 ;
        RECT 47.338 62.969 54.116 63.027 ;
        RECT 47.292 63.015 54.07 63.073 ;
        RECT 47.246 63.061 54.024 63.119 ;
        RECT 47.2 63.107 53.978 63.165 ;
        RECT 47.154 63.153 53.932 63.211 ;
        RECT 47.108 63.199 53.886 63.257 ;
        RECT 47.062 63.245 53.84 63.303 ;
        RECT 47.016 63.291 53.794 63.349 ;
        RECT 46.97 63.337 53.748 63.395 ;
        RECT 46.924 63.383 53.702 63.441 ;
        RECT 46.878 63.429 53.656 63.487 ;
        RECT 46.832 63.475 53.61 63.533 ;
        RECT 46.786 63.521 53.564 63.579 ;
        RECT 46.74 63.567 53.518 63.625 ;
        RECT 46.694 63.613 53.472 63.671 ;
        RECT 46.648 63.659 53.426 63.717 ;
        RECT 46.602 63.705 53.38 63.763 ;
        RECT 46.556 63.751 53.334 63.809 ;
        RECT 46.51 63.797 53.288 63.855 ;
        RECT 46.464 63.843 53.242 63.901 ;
        RECT 46.418 63.889 53.196 63.947 ;
        RECT 46.372 63.935 53.15 63.993 ;
        RECT 46.326 63.981 53.104 64.039 ;
        RECT 46.28 64.027 53.058 64.085 ;
        RECT 46.234 64.073 53.012 64.131 ;
        RECT 46.188 64.119 52.966 64.177 ;
        RECT 46.142 64.165 52.92 64.223 ;
        RECT 46.096 64.211 52.874 64.269 ;
        RECT 46.05 64.257 52.828 64.315 ;
        RECT 46.004 64.303 52.782 64.361 ;
        RECT 45.958 64.349 52.736 64.407 ;
        RECT 45.912 64.395 52.69 64.453 ;
        RECT 45.866 64.441 52.644 64.499 ;
        RECT 45.82 64.487 52.598 64.545 ;
        RECT 45.774 64.533 52.552 64.591 ;
        RECT 45.728 64.579 52.506 64.637 ;
        RECT 45.682 64.625 52.46 64.683 ;
        RECT 45.636 64.671 52.414 64.729 ;
        RECT 45.59 64.717 52.368 64.775 ;
        RECT 45.544 64.763 52.322 64.821 ;
        RECT 45.498 64.809 52.276 64.867 ;
        RECT 45.452 64.855 52.23 64.913 ;
        RECT 45.406 64.901 52.184 64.959 ;
        RECT 45.36 64.947 52.138 65.005 ;
        RECT 45.314 64.993 52.092 65.051 ;
        RECT 45.268 65.039 52.046 65.097 ;
        RECT 45.222 65.085 52 65.143 ;
        RECT 45.176 65.131 51.954 65.189 ;
        RECT 45.13 65.177 51.908 65.235 ;
        RECT 45.084 65.223 51.862 65.281 ;
        RECT 45.038 65.269 51.816 65.327 ;
        RECT 44.992 65.315 51.77 65.373 ;
        RECT 44.946 65.361 51.724 65.419 ;
        RECT 44.9 65.407 51.678 65.465 ;
        RECT 44.854 65.453 51.632 65.511 ;
        RECT 44.808 65.499 51.586 65.557 ;
        RECT 44.762 65.545 51.54 65.603 ;
        RECT 44.716 65.591 51.494 65.649 ;
        RECT 44.67 65.637 51.448 65.695 ;
        RECT 44.624 65.683 51.402 65.741 ;
        RECT 44.578 65.729 51.356 65.787 ;
        RECT 44.532 65.775 51.31 65.833 ;
        RECT 44.486 65.821 51.264 65.879 ;
        RECT 44.44 65.867 51.218 65.925 ;
        RECT 44.394 65.913 51.172 65.971 ;
        RECT 44.348 65.959 51.126 66.017 ;
        RECT 44.302 66.005 51.08 66.063 ;
        RECT 44.256 66.051 51.034 66.109 ;
        RECT 44.21 66.097 50.988 66.155 ;
        RECT 44.164 66.143 50.942 66.201 ;
        RECT 44.118 66.189 50.896 66.247 ;
        RECT 44.072 66.235 50.85 66.293 ;
        RECT 44.026 66.281 50.804 66.339 ;
        RECT 43.98 66.327 50.758 66.385 ;
        RECT 43.934 66.373 50.712 66.431 ;
        RECT 43.888 66.419 50.666 66.477 ;
        RECT 43.842 66.465 50.62 66.523 ;
        RECT 43.796 66.511 50.574 66.569 ;
        RECT 43.75 66.557 50.528 66.615 ;
        RECT 43.704 66.603 50.482 66.661 ;
        RECT 43.658 66.649 50.436 66.707 ;
        RECT 43.612 66.695 50.39 66.753 ;
        RECT 43.566 66.741 50.344 66.799 ;
        RECT 43.52 66.787 50.298 66.845 ;
        RECT 43.474 66.833 50.252 66.891 ;
        RECT 43.428 66.879 50.206 66.937 ;
        RECT 43.382 66.925 50.16 66.983 ;
        RECT 43.336 66.971 50.114 67.029 ;
        RECT 43.29 67.017 50.068 67.075 ;
        RECT 43.244 67.063 50.022 67.121 ;
        RECT 43.198 67.109 49.976 67.167 ;
        RECT 43.152 67.155 49.93 67.213 ;
        RECT 43.106 67.201 49.884 67.259 ;
        RECT 43.06 67.247 49.838 67.305 ;
        RECT 43.014 67.293 49.792 67.351 ;
        RECT 42.968 67.339 49.746 67.397 ;
        RECT 42.922 67.385 49.7 67.443 ;
        RECT 42.876 67.431 49.654 67.489 ;
        RECT 42.83 67.477 49.608 67.535 ;
        RECT 42.784 67.523 49.562 67.581 ;
        RECT 42.738 67.569 49.516 67.627 ;
        RECT 42.692 67.615 49.47 67.673 ;
        RECT 42.646 67.661 49.424 67.719 ;
        RECT 42.6 67.707 49.378 67.765 ;
        RECT 42.6 67.707 49.332 67.811 ;
        RECT 42.6 67.707 49.286 67.857 ;
        RECT 42.6 67.707 49.24 67.903 ;
        RECT 42.6 67.707 49.194 67.949 ;
        RECT 42.6 67.707 49.148 67.995 ;
        RECT 42.6 67.707 49.102 68.041 ;
        RECT 42.6 67.707 49.056 68.087 ;
        RECT 42.6 67.707 49.01 68.133 ;
        RECT 42.6 67.707 48.964 68.179 ;
        RECT 42.6 67.707 48.918 68.225 ;
        RECT 42.6 67.707 48.872 68.271 ;
        RECT 42.6 67.707 48.826 68.317 ;
        RECT 42.6 67.707 48.78 68.363 ;
        RECT 42.6 67.707 48.734 68.409 ;
        RECT 42.6 67.707 48.688 68.455 ;
        RECT 42.6 67.707 48.642 68.501 ;
        RECT 42.6 67.707 48.596 68.547 ;
        RECT 42.6 67.707 48.55 68.593 ;
        RECT 42.6 67.707 48.504 68.639 ;
        RECT 42.6 67.707 48.458 68.685 ;
        RECT 42.6 67.707 48.412 68.731 ;
        RECT 42.6 67.707 48.366 68.777 ;
        RECT 42.6 67.707 48.32 68.823 ;
        RECT 42.6 67.707 48.274 68.869 ;
        RECT 42.6 67.707 48.228 68.915 ;
        RECT 42.6 67.707 48.182 68.961 ;
        RECT 42.6 67.707 48.136 69.007 ;
        RECT 42.6 67.707 48.09 69.053 ;
        RECT 42.6 67.707 48.044 69.099 ;
        RECT 42.6 67.707 47.998 69.145 ;
        RECT 42.6 67.707 47.952 69.191 ;
        RECT 42.6 67.707 47.906 69.237 ;
        RECT 42.6 67.707 47.86 69.283 ;
        RECT 42.6 67.707 47.814 69.329 ;
        RECT 42.6 67.707 47.768 69.375 ;
        RECT 42.6 67.707 47.722 69.421 ;
        RECT 42.6 67.707 47.676 69.467 ;
        RECT 42.6 67.707 47.63 69.513 ;
        RECT 42.6 67.707 47.584 69.559 ;
        RECT 42.6 67.707 47.538 69.605 ;
        RECT 42.6 67.707 47.492 69.651 ;
        RECT 42.6 67.707 47.446 69.697 ;
        RECT 42.6 67.707 47.4 80 ;
    END
    PORT
      LAYER QB ;
        RECT 32.076 51.921 38.838 51.995 ;
        RECT 32.03 51.967 38.792 52.041 ;
        RECT 31.984 52.013 38.746 52.087 ;
        RECT 31.938 52.059 38.7 52.133 ;
        RECT 31.892 52.105 38.654 52.179 ;
        RECT 31.846 52.151 38.608 52.225 ;
        RECT 31.8 52.197 38.562 52.271 ;
        RECT 31.754 52.243 38.516 52.317 ;
        RECT 31.708 52.289 38.47 52.363 ;
        RECT 31.662 52.335 38.424 52.409 ;
        RECT 31.616 52.381 38.378 52.455 ;
        RECT 31.57 52.427 38.332 52.501 ;
        RECT 31.524 52.473 38.286 52.547 ;
        RECT 31.478 52.519 38.24 52.593 ;
        RECT 31.432 52.565 38.194 52.639 ;
        RECT 31.386 52.611 38.148 52.685 ;
        RECT 31.34 52.657 38.102 52.731 ;
        RECT 31.294 52.703 38.056 52.777 ;
        RECT 31.248 52.749 38.01 52.823 ;
        RECT 31.202 52.795 37.964 52.869 ;
        RECT 31.156 52.841 37.918 52.915 ;
        RECT 31.11 52.887 37.872 52.961 ;
        RECT 31.064 52.933 37.826 53.007 ;
        RECT 31.018 52.979 37.78 53.053 ;
        RECT 30.972 53.025 37.734 53.099 ;
        RECT 30.926 53.071 37.688 53.145 ;
        RECT 30.88 53.117 37.642 53.191 ;
        RECT 30.834 53.163 37.596 53.237 ;
        RECT 30.788 53.209 37.55 53.283 ;
        RECT 30.742 53.255 37.504 53.329 ;
        RECT 30.696 53.301 37.458 53.375 ;
        RECT 30.65 53.347 37.412 53.421 ;
        RECT 30.604 53.393 37.366 53.467 ;
        RECT 30.558 53.439 37.32 53.513 ;
        RECT 30.512 53.485 37.274 53.559 ;
        RECT 30.466 53.531 37.228 53.605 ;
        RECT 30.42 53.577 37.182 53.651 ;
        RECT 30.374 53.623 37.136 53.697 ;
        RECT 30.328 53.669 37.09 53.743 ;
        RECT 30.282 53.715 37.044 53.789 ;
        RECT 30.236 53.761 36.998 53.835 ;
        RECT 30.19 53.807 36.952 53.881 ;
        RECT 30.144 53.853 36.906 53.927 ;
        RECT 30.098 53.899 36.86 53.973 ;
        RECT 30.052 53.945 36.814 54.019 ;
        RECT 30.006 53.991 36.768 54.065 ;
        RECT 29.96 54.037 36.722 54.111 ;
        RECT 29.914 54.083 36.676 54.157 ;
        RECT 29.868 54.129 36.63 54.203 ;
        RECT 29.822 54.175 36.584 54.249 ;
        RECT 29.776 54.221 36.538 54.295 ;
        RECT 29.73 54.267 36.492 54.341 ;
        RECT 29.684 54.313 36.446 54.387 ;
        RECT 29.638 54.359 36.4 54.433 ;
        RECT 29.592 54.405 36.354 54.479 ;
        RECT 29.546 54.451 36.308 54.525 ;
        RECT 29.5 54.497 36.262 54.571 ;
        RECT 29.454 54.543 36.216 54.617 ;
        RECT 29.408 54.589 36.17 54.663 ;
        RECT 29.362 54.635 36.124 54.709 ;
        RECT 29.316 54.681 36.078 54.755 ;
        RECT 29.27 54.727 36.032 54.801 ;
        RECT 29.224 54.773 35.986 54.847 ;
        RECT 29.178 54.819 35.94 54.893 ;
        RECT 29.132 54.865 35.894 54.939 ;
        RECT 29.086 54.911 35.848 54.985 ;
        RECT 29.04 54.957 35.802 55.031 ;
        RECT 28.994 55.003 35.756 55.077 ;
        RECT 28.948 55.049 35.71 55.123 ;
        RECT 28.902 55.095 35.664 55.169 ;
        RECT 28.856 55.141 35.618 55.215 ;
        RECT 28.81 55.187 35.572 55.261 ;
        RECT 28.764 55.233 35.526 55.307 ;
        RECT 28.718 55.279 35.48 55.353 ;
        RECT 28.672 55.325 35.434 55.399 ;
        RECT 28.626 55.371 35.388 55.445 ;
        RECT 28.58 55.417 35.342 55.491 ;
        RECT 28.534 55.463 35.296 55.537 ;
        RECT 28.488 55.509 35.25 55.583 ;
        RECT 28.442 55.555 35.204 55.629 ;
        RECT 28.396 55.601 35.158 55.675 ;
        RECT 28.35 55.647 35.112 55.721 ;
        RECT 28.304 55.693 35.066 55.767 ;
        RECT 28.258 55.739 35.02 55.813 ;
        RECT 28.212 55.785 34.974 55.859 ;
        RECT 28.166 55.831 34.928 55.905 ;
        RECT 28.12 55.877 34.882 55.951 ;
        RECT 28.074 55.923 34.836 55.997 ;
        RECT 28.028 55.969 34.79 56.043 ;
        RECT 27.982 56.015 34.744 56.089 ;
        RECT 27.936 56.061 34.698 56.135 ;
        RECT 27.89 56.107 34.652 56.181 ;
        RECT 27.844 56.153 34.606 56.227 ;
        RECT 27.798 56.199 34.56 56.273 ;
        RECT 27.752 56.245 34.514 56.319 ;
        RECT 27.706 56.291 34.468 56.365 ;
        RECT 27.66 56.337 34.422 56.411 ;
        RECT 27.614 56.383 34.376 56.457 ;
        RECT 27.568 56.429 34.33 56.503 ;
        RECT 27.522 56.475 34.284 56.549 ;
        RECT 27.476 56.521 34.238 56.595 ;
        RECT 27.43 56.567 34.192 56.641 ;
        RECT 27.384 56.613 34.146 56.687 ;
        RECT 27.338 56.659 34.1 56.733 ;
        RECT 27.292 56.705 34.054 56.779 ;
        RECT 27.246 56.751 34.008 56.825 ;
        RECT 27.2 56.797 33.962 56.871 ;
        RECT 27.154 56.843 33.916 56.917 ;
        RECT 27.108 56.889 33.87 56.963 ;
        RECT 27.062 56.935 33.824 57.009 ;
        RECT 27.016 56.981 33.778 57.055 ;
        RECT 26.97 57.027 33.732 57.101 ;
        RECT 26.924 57.073 33.686 57.147 ;
        RECT 26.878 57.119 33.64 57.193 ;
        RECT 26.832 57.165 33.594 57.239 ;
        RECT 26.786 57.211 33.548 57.285 ;
        RECT 26.74 57.257 33.502 57.331 ;
        RECT 26.694 57.303 33.456 57.377 ;
        RECT 26.648 57.349 33.41 57.423 ;
        RECT 26.602 57.395 33.364 57.469 ;
        RECT 26.556 57.441 33.318 57.515 ;
        RECT 26.51 57.487 33.272 57.561 ;
        RECT 26.464 57.533 33.226 57.607 ;
        RECT 26.418 57.579 33.18 57.653 ;
        RECT 26.372 57.625 33.134 57.699 ;
        RECT 26.326 57.671 33.088 57.745 ;
        RECT 26.28 57.717 33.042 57.791 ;
        RECT 26.234 57.763 32.996 57.837 ;
        RECT 26.188 57.809 32.95 57.883 ;
        RECT 26.142 57.855 32.904 57.929 ;
        RECT 26.096 57.901 32.858 57.975 ;
        RECT 26.05 57.947 32.812 58.021 ;
        RECT 26.004 57.993 32.766 58.067 ;
        RECT 25.958 58.039 32.72 58.113 ;
        RECT 25.912 58.085 32.674 58.159 ;
        RECT 25.866 58.131 32.628 58.205 ;
        RECT 25.82 58.177 32.582 58.251 ;
        RECT 25.774 58.223 32.536 58.297 ;
        RECT 25.728 58.269 32.49 58.343 ;
        RECT 25.682 58.315 32.444 58.389 ;
        RECT 25.636 58.361 32.398 58.435 ;
        RECT 25.59 58.407 32.352 58.481 ;
        RECT 25.544 58.453 32.306 58.527 ;
        RECT 25.498 58.499 32.26 58.573 ;
        RECT 25.452 58.545 32.214 58.619 ;
        RECT 25.406 58.591 32.168 58.665 ;
        RECT 25.36 58.637 32.122 58.711 ;
        RECT 25.314 58.683 32.076 58.757 ;
        RECT 25.268 58.729 32.03 58.803 ;
        RECT 25.222 58.775 31.984 58.849 ;
        RECT 25.176 58.821 31.938 58.895 ;
        RECT 25.13 58.867 31.892 58.941 ;
        RECT 25.084 58.913 31.846 58.987 ;
        RECT 25.038 58.959 31.8 59.033 ;
        RECT 24.992 59.005 31.754 59.079 ;
        RECT 24.946 59.051 31.708 59.125 ;
        RECT 24.9 59.097 31.662 59.171 ;
        RECT 24.854 59.143 31.616 59.217 ;
        RECT 24.808 59.189 31.57 59.263 ;
        RECT 24.762 59.235 31.524 59.309 ;
        RECT 24.716 59.281 31.478 59.355 ;
        RECT 24.67 59.327 31.432 59.401 ;
        RECT 24.624 59.373 31.386 59.447 ;
        RECT 24.578 59.419 31.34 59.493 ;
        RECT 24.532 59.465 31.294 59.539 ;
        RECT 24.486 59.511 31.248 59.585 ;
        RECT 24.44 59.557 31.202 59.631 ;
        RECT 24.394 59.603 31.156 59.677 ;
        RECT 24.348 59.649 31.11 59.723 ;
        RECT 24.302 59.695 31.064 59.769 ;
        RECT 24.256 59.741 31.018 59.815 ;
        RECT 24.21 59.787 30.972 59.861 ;
        RECT 24.164 59.833 30.926 59.907 ;
        RECT 24.118 59.879 30.88 59.953 ;
        RECT 24.072 59.925 30.834 59.999 ;
        RECT 24.026 59.971 30.788 60.045 ;
        RECT 23.98 60.017 30.742 60.091 ;
        RECT 23.934 60.063 30.696 60.137 ;
        RECT 23.888 60.109 30.65 60.183 ;
        RECT 23.842 60.155 30.604 60.229 ;
        RECT 23.796 60.201 30.558 60.275 ;
        RECT 23.75 60.247 30.512 60.321 ;
        RECT 23.704 60.293 30.466 60.367 ;
        RECT 23.658 60.339 30.42 60.413 ;
        RECT 23.612 60.385 30.374 60.459 ;
        RECT 23.566 60.431 30.328 60.505 ;
        RECT 23.52 60.477 30.282 60.551 ;
        RECT 23.474 60.523 30.236 60.597 ;
        RECT 23.428 60.569 30.19 60.643 ;
        RECT 23.382 60.615 30.144 60.689 ;
        RECT 23.336 60.661 30.098 60.735 ;
        RECT 23.29 60.707 30.052 60.781 ;
        RECT 23.244 60.753 30.006 60.827 ;
        RECT 23.198 60.799 29.96 60.873 ;
        RECT 23.152 60.845 29.914 60.919 ;
        RECT 23.106 60.891 29.868 60.965 ;
        RECT 23.06 60.937 29.822 61.011 ;
        RECT 23.014 60.983 29.776 61.057 ;
        RECT 22.968 61.029 29.73 61.103 ;
        RECT 22.922 61.075 29.684 61.149 ;
        RECT 22.876 61.121 29.638 61.195 ;
        RECT 22.83 61.167 29.592 61.241 ;
        RECT 22.784 61.213 29.546 61.287 ;
        RECT 22.738 61.259 29.5 61.333 ;
        RECT 22.692 61.305 29.454 61.379 ;
        RECT 22.646 61.351 29.408 61.425 ;
        RECT 22.584 61.428 29.362 61.471 ;
        RECT 22.6 61.397 29.362 61.471 ;
        RECT 22.538 61.459 29.316 61.517 ;
        RECT 22.492 61.505 29.27 61.563 ;
        RECT 22.446 61.551 29.224 61.609 ;
        RECT 22.4 61.597 29.178 61.655 ;
        RECT 22.354 61.643 29.132 61.701 ;
        RECT 22.308 61.689 29.086 61.747 ;
        RECT 22.262 61.735 29.04 61.793 ;
        RECT 22.216 61.781 28.994 61.839 ;
        RECT 22.17 61.827 28.948 61.885 ;
        RECT 22.124 61.873 28.902 61.931 ;
        RECT 22.078 61.919 28.856 61.977 ;
        RECT 22.032 61.965 28.81 62.023 ;
        RECT 21.986 62.011 28.764 62.069 ;
        RECT 21.94 62.057 28.718 62.115 ;
        RECT 21.894 62.103 28.672 62.161 ;
        RECT 21.848 62.149 28.626 62.207 ;
        RECT 21.802 62.195 28.58 62.253 ;
        RECT 21.756 62.241 28.534 62.299 ;
        RECT 21.71 62.287 28.488 62.345 ;
        RECT 21.664 62.333 28.442 62.391 ;
        RECT 21.618 62.379 28.396 62.437 ;
        RECT 21.572 62.425 28.35 62.483 ;
        RECT 21.526 62.471 28.304 62.529 ;
        RECT 21.48 62.517 28.258 62.575 ;
        RECT 21.434 62.563 28.212 62.621 ;
        RECT 21.388 62.609 28.166 62.667 ;
        RECT 21.342 62.655 28.12 62.713 ;
        RECT 21.296 62.701 28.074 62.759 ;
        RECT 21.25 62.747 28.028 62.805 ;
        RECT 21.204 62.793 27.982 62.851 ;
        RECT 21.158 62.839 27.936 62.897 ;
        RECT 21.112 62.885 27.89 62.943 ;
        RECT 21.066 62.931 27.844 62.989 ;
        RECT 21.02 62.977 27.798 63.035 ;
        RECT 20.974 63.023 27.752 63.081 ;
        RECT 20.928 63.069 27.706 63.127 ;
        RECT 20.882 63.115 27.66 63.173 ;
        RECT 20.836 63.161 27.614 63.219 ;
        RECT 20.79 63.207 27.568 63.265 ;
        RECT 20.744 63.253 27.522 63.311 ;
        RECT 20.698 63.299 27.476 63.357 ;
        RECT 20.652 63.345 27.43 63.403 ;
        RECT 20.606 63.391 27.384 63.449 ;
        RECT 20.56 63.437 27.338 63.495 ;
        RECT 20.514 63.483 27.292 63.541 ;
        RECT 20.468 63.529 27.246 63.587 ;
        RECT 20.422 63.575 27.2 63.633 ;
        RECT 20.376 63.621 27.154 63.679 ;
        RECT 20.33 63.667 27.108 63.725 ;
        RECT 20.284 63.713 27.062 63.771 ;
        RECT 20.238 63.759 27.016 63.817 ;
        RECT 20.192 63.805 26.97 63.863 ;
        RECT 20.146 63.851 26.924 63.909 ;
        RECT 20.1 63.897 26.878 63.955 ;
        RECT 20.054 63.943 26.832 64.001 ;
        RECT 20.008 63.989 26.786 64.047 ;
        RECT 19.962 64.035 26.74 64.093 ;
        RECT 19.916 64.081 26.694 64.139 ;
        RECT 19.87 64.127 26.648 64.185 ;
        RECT 19.824 64.173 26.602 64.231 ;
        RECT 19.778 64.219 26.556 64.277 ;
        RECT 19.732 64.265 26.51 64.323 ;
        RECT 19.686 64.311 26.464 64.369 ;
        RECT 19.64 64.357 26.418 64.415 ;
        RECT 19.594 64.403 26.372 64.461 ;
        RECT 19.548 64.449 26.326 64.507 ;
        RECT 19.502 64.495 26.28 64.553 ;
        RECT 19.456 64.541 26.234 64.599 ;
        RECT 19.41 64.587 26.188 64.645 ;
        RECT 19.364 64.633 26.142 64.691 ;
        RECT 19.318 64.679 26.096 64.737 ;
        RECT 19.272 64.725 26.05 64.783 ;
        RECT 19.226 64.771 26.004 64.829 ;
        RECT 19.18 64.817 25.958 64.875 ;
        RECT 19.134 64.863 25.912 64.921 ;
        RECT 19.088 64.909 25.866 64.967 ;
        RECT 19.042 64.955 25.82 65.013 ;
        RECT 18.996 65.001 25.774 65.059 ;
        RECT 18.95 65.047 25.728 65.105 ;
        RECT 18.904 65.093 25.682 65.151 ;
        RECT 18.858 65.139 25.636 65.197 ;
        RECT 18.812 65.185 25.59 65.243 ;
        RECT 18.766 65.231 25.544 65.289 ;
        RECT 18.72 65.277 25.498 65.335 ;
        RECT 18.674 65.323 25.452 65.381 ;
        RECT 18.628 65.369 25.406 65.427 ;
        RECT 18.582 65.415 25.36 65.473 ;
        RECT 18.536 65.461 25.314 65.519 ;
        RECT 18.49 65.507 25.268 65.565 ;
        RECT 18.444 65.553 25.222 65.611 ;
        RECT 18.398 65.599 25.176 65.657 ;
        RECT 18.352 65.645 25.13 65.703 ;
        RECT 18.306 65.691 25.084 65.749 ;
        RECT 18.26 65.737 25.038 65.795 ;
        RECT 18.214 65.783 24.992 65.841 ;
        RECT 18.168 65.829 24.946 65.887 ;
        RECT 18.122 65.875 24.9 65.933 ;
        RECT 18.076 65.921 24.854 65.979 ;
        RECT 18.03 65.967 24.808 66.025 ;
        RECT 17.984 66.013 24.762 66.071 ;
        RECT 17.938 66.059 24.716 66.117 ;
        RECT 17.892 66.105 24.67 66.163 ;
        RECT 17.846 66.151 24.624 66.209 ;
        RECT 17.8 66.197 24.578 66.255 ;
        RECT 17.8 66.197 24.532 66.301 ;
        RECT 17.8 66.197 24.486 66.347 ;
        RECT 17.8 66.197 24.44 66.393 ;
        RECT 17.8 66.197 24.394 66.439 ;
        RECT 17.8 66.197 24.348 66.485 ;
        RECT 17.8 66.197 24.302 66.531 ;
        RECT 17.8 66.197 24.256 66.577 ;
        RECT 17.8 66.197 24.21 66.623 ;
        RECT 17.8 66.197 24.164 66.669 ;
        RECT 17.8 66.197 24.118 66.715 ;
        RECT 17.8 66.197 24.072 66.761 ;
        RECT 17.8 66.197 24.026 66.807 ;
        RECT 17.8 66.197 23.98 66.853 ;
        RECT 17.8 66.197 23.934 66.899 ;
        RECT 17.8 66.197 23.888 66.945 ;
        RECT 17.8 66.197 23.842 66.991 ;
        RECT 17.8 66.197 23.796 67.037 ;
        RECT 17.8 66.197 23.75 67.083 ;
        RECT 17.8 66.197 23.704 67.129 ;
        RECT 17.8 66.197 23.658 67.175 ;
        RECT 17.8 66.197 23.612 67.221 ;
        RECT 17.8 66.197 23.566 67.267 ;
        RECT 17.8 66.197 23.52 67.313 ;
        RECT 17.8 66.197 23.474 67.359 ;
        RECT 17.8 66.197 23.428 67.405 ;
        RECT 17.8 66.197 23.382 67.451 ;
        RECT 17.8 66.197 23.336 67.497 ;
        RECT 17.8 66.197 23.29 67.543 ;
        RECT 17.8 66.197 23.244 67.589 ;
        RECT 17.8 66.197 23.198 67.635 ;
        RECT 17.8 66.197 23.152 67.681 ;
        RECT 17.8 66.197 23.106 67.727 ;
        RECT 17.8 66.197 23.06 67.773 ;
        RECT 17.8 66.197 23.014 67.819 ;
        RECT 17.8 66.197 22.968 67.865 ;
        RECT 17.8 66.197 22.922 67.911 ;
        RECT 17.8 66.197 22.876 67.957 ;
        RECT 17.8 66.197 22.83 68.003 ;
        RECT 17.8 66.197 22.784 68.049 ;
        RECT 17.8 66.197 22.738 68.095 ;
        RECT 17.8 66.197 22.692 68.141 ;
        RECT 17.8 66.197 22.646 68.187 ;
        RECT 17.8 66.197 22.6 80 ;
        RECT 66.22 17.8 80 22.6 ;
        RECT 61.424 22.573 68.21 22.606 ;
        RECT 59.446 24.551 66.22 24.596 ;
        RECT 59.492 24.505 66.266 24.567 ;
        RECT 66.208 17.806 66.22 24.596 ;
        RECT 59.538 24.459 66.312 24.521 ;
        RECT 66.162 17.835 66.208 24.625 ;
        RECT 59.4 24.597 66.162 24.671 ;
        RECT 59.584 24.413 66.358 24.475 ;
        RECT 66.116 17.881 66.162 24.671 ;
        RECT 59.354 24.643 66.116 24.717 ;
        RECT 59.63 24.367 66.404 24.429 ;
        RECT 66.07 17.927 66.116 24.717 ;
        RECT 59.308 24.689 66.07 24.763 ;
        RECT 59.676 24.321 66.45 24.383 ;
        RECT 66.024 17.973 66.07 24.763 ;
        RECT 59.262 24.735 66.024 24.809 ;
        RECT 59.722 24.275 66.496 24.337 ;
        RECT 65.978 18.019 66.024 24.809 ;
        RECT 59.216 24.781 65.978 24.855 ;
        RECT 59.768 24.229 66.542 24.291 ;
        RECT 65.932 18.065 65.978 24.855 ;
        RECT 59.17 24.827 65.932 24.901 ;
        RECT 59.814 24.183 66.588 24.245 ;
        RECT 65.886 18.111 65.932 24.901 ;
        RECT 59.124 24.873 65.886 24.947 ;
        RECT 59.86 24.137 66.634 24.199 ;
        RECT 65.84 18.157 65.886 24.947 ;
        RECT 59.078 24.919 65.84 24.993 ;
        RECT 59.906 24.091 66.68 24.153 ;
        RECT 65.794 18.203 65.84 24.993 ;
        RECT 59.032 24.965 65.794 25.039 ;
        RECT 59.952 24.045 66.726 24.107 ;
        RECT 65.748 18.249 65.794 25.039 ;
        RECT 58.986 25.011 65.748 25.085 ;
        RECT 59.998 23.999 66.772 24.061 ;
        RECT 65.702 18.295 65.748 25.085 ;
        RECT 58.94 25.057 65.702 25.131 ;
        RECT 60.044 23.953 66.818 24.015 ;
        RECT 65.656 18.341 65.702 25.131 ;
        RECT 58.894 25.103 65.656 25.177 ;
        RECT 60.09 23.907 66.864 23.969 ;
        RECT 65.61 18.387 65.656 25.177 ;
        RECT 58.848 25.149 65.61 25.223 ;
        RECT 60.136 23.861 66.91 23.923 ;
        RECT 65.564 18.433 65.61 25.223 ;
        RECT 58.802 25.195 65.564 25.269 ;
        RECT 60.182 23.815 66.956 23.877 ;
        RECT 65.518 18.479 65.564 25.269 ;
        RECT 58.756 25.241 65.518 25.315 ;
        RECT 60.228 23.769 67.002 23.831 ;
        RECT 65.472 18.525 65.518 25.315 ;
        RECT 58.71 25.287 65.472 25.361 ;
        RECT 60.274 23.723 67.048 23.785 ;
        RECT 65.426 18.571 65.472 25.361 ;
        RECT 58.664 25.333 65.426 25.407 ;
        RECT 60.32 23.677 67.094 23.739 ;
        RECT 65.38 18.617 65.426 25.407 ;
        RECT 58.618 25.379 65.38 25.453 ;
        RECT 60.366 23.631 67.14 23.693 ;
        RECT 65.334 18.663 65.38 25.453 ;
        RECT 58.572 25.425 65.334 25.499 ;
        RECT 60.412 23.585 67.186 23.647 ;
        RECT 65.288 18.709 65.334 25.499 ;
        RECT 58.526 25.471 65.288 25.545 ;
        RECT 60.458 23.539 67.232 23.601 ;
        RECT 65.242 18.755 65.288 25.545 ;
        RECT 58.48 25.517 65.242 25.591 ;
        RECT 60.504 23.493 67.278 23.555 ;
        RECT 65.196 18.801 65.242 25.591 ;
        RECT 58.434 25.563 65.196 25.637 ;
        RECT 60.55 23.447 67.324 23.509 ;
        RECT 65.15 18.847 65.196 25.637 ;
        RECT 58.388 25.609 65.15 25.683 ;
        RECT 60.596 23.401 67.37 23.463 ;
        RECT 65.104 18.893 65.15 25.683 ;
        RECT 58.342 25.655 65.104 25.729 ;
        RECT 60.642 23.355 67.416 23.417 ;
        RECT 65.058 18.939 65.104 25.729 ;
        RECT 58.296 25.701 65.058 25.775 ;
        RECT 60.688 23.309 67.462 23.371 ;
        RECT 65.012 18.985 65.058 25.775 ;
        RECT 58.25 25.747 65.012 25.821 ;
        RECT 60.734 23.263 67.508 23.325 ;
        RECT 64.966 19.031 65.012 25.821 ;
        RECT 58.204 25.793 64.966 25.867 ;
        RECT 60.78 23.217 67.554 23.279 ;
        RECT 64.92 19.077 64.966 25.867 ;
        RECT 58.158 25.839 64.92 25.913 ;
        RECT 60.826 23.171 67.6 23.233 ;
        RECT 64.874 19.123 64.92 25.913 ;
        RECT 58.112 25.885 64.874 25.959 ;
        RECT 60.872 23.125 67.646 23.187 ;
        RECT 64.828 19.169 64.874 25.959 ;
        RECT 58.066 25.931 64.828 26.005 ;
        RECT 60.918 23.079 67.692 23.141 ;
        RECT 64.782 19.215 64.828 26.005 ;
        RECT 58.02 25.977 64.782 26.051 ;
        RECT 60.964 23.033 67.738 23.095 ;
        RECT 64.736 19.261 64.782 26.051 ;
        RECT 57.974 26.023 64.736 26.097 ;
        RECT 61.01 22.987 67.784 23.049 ;
        RECT 64.69 19.307 64.736 26.097 ;
        RECT 57.928 26.069 64.69 26.143 ;
        RECT 61.056 22.941 67.83 23.003 ;
        RECT 64.644 19.353 64.69 26.143 ;
        RECT 57.882 26.115 64.644 26.189 ;
        RECT 61.102 22.895 67.876 22.957 ;
        RECT 64.598 19.399 64.644 26.189 ;
        RECT 57.836 26.161 64.598 26.235 ;
        RECT 61.148 22.849 67.922 22.911 ;
        RECT 64.552 19.445 64.598 26.235 ;
        RECT 57.79 26.207 64.552 26.281 ;
        RECT 61.194 22.803 67.968 22.865 ;
        RECT 64.506 19.491 64.552 26.281 ;
        RECT 57.744 26.253 64.506 26.327 ;
        RECT 61.24 22.757 68.014 22.819 ;
        RECT 64.46 19.537 64.506 26.327 ;
        RECT 57.698 26.299 64.46 26.373 ;
        RECT 61.286 22.711 68.06 22.773 ;
        RECT 64.414 19.583 64.46 26.373 ;
        RECT 57.652 26.345 64.414 26.419 ;
        RECT 61.332 22.665 68.106 22.727 ;
        RECT 64.368 19.629 64.414 26.419 ;
        RECT 57.606 26.391 64.368 26.465 ;
        RECT 61.378 22.619 68.152 22.681 ;
        RECT 64.322 19.675 64.368 26.465 ;
        RECT 57.56 26.437 64.322 26.511 ;
        RECT 61.424 22.573 68.198 22.635 ;
        RECT 64.276 19.721 64.322 26.511 ;
        RECT 57.514 26.483 64.276 26.557 ;
        RECT 61.47 22.527 80 22.6 ;
        RECT 64.23 19.767 64.276 26.557 ;
        RECT 57.468 26.529 64.23 26.603 ;
        RECT 61.516 22.481 80 22.6 ;
        RECT 64.184 19.813 64.23 26.603 ;
        RECT 57.422 26.575 64.184 26.649 ;
        RECT 61.562 22.435 80 22.6 ;
        RECT 64.138 19.859 64.184 26.649 ;
        RECT 57.376 26.621 64.138 26.695 ;
        RECT 61.608 22.389 80 22.6 ;
        RECT 64.092 19.905 64.138 26.695 ;
        RECT 57.33 26.667 64.092 26.741 ;
        RECT 61.654 22.343 80 22.6 ;
        RECT 64.046 19.951 64.092 26.741 ;
        RECT 57.284 26.713 64.046 26.787 ;
        RECT 61.7 22.297 80 22.6 ;
        RECT 64 19.997 64.046 26.787 ;
        RECT 57.238 26.759 64 26.833 ;
        RECT 61.746 22.251 80 22.6 ;
        RECT 63.954 20.043 64 26.833 ;
        RECT 57.192 26.805 63.954 26.879 ;
        RECT 61.792 22.205 80 22.6 ;
        RECT 63.908 20.089 63.954 26.879 ;
        RECT 57.146 26.851 63.908 26.925 ;
        RECT 61.838 22.159 80 22.6 ;
        RECT 63.862 20.135 63.908 26.925 ;
        RECT 57.1 26.897 63.862 26.971 ;
        RECT 61.884 22.113 80 22.6 ;
        RECT 63.816 20.181 63.862 26.971 ;
        RECT 57.054 26.943 63.816 27.017 ;
        RECT 61.93 22.067 80 22.6 ;
        RECT 63.77 20.227 63.816 27.017 ;
        RECT 57.008 26.989 63.77 27.063 ;
        RECT 61.976 22.021 80 22.6 ;
        RECT 63.724 20.273 63.77 27.063 ;
        RECT 56.962 27.035 63.724 27.109 ;
        RECT 62.022 21.975 80 22.6 ;
        RECT 63.678 20.319 63.724 27.109 ;
        RECT 56.916 27.081 63.678 27.155 ;
        RECT 62.068 21.929 80 22.6 ;
        RECT 63.632 20.365 63.678 27.155 ;
        RECT 56.87 27.127 63.632 27.201 ;
        RECT 62.114 21.883 80 22.6 ;
        RECT 63.586 20.411 63.632 27.201 ;
        RECT 56.824 27.173 63.586 27.247 ;
        RECT 62.16 21.837 80 22.6 ;
        RECT 63.54 20.457 63.586 27.247 ;
        RECT 56.778 27.219 63.54 27.293 ;
        RECT 62.206 21.791 80 22.6 ;
        RECT 63.494 20.503 63.54 27.293 ;
        RECT 56.732 27.265 63.494 27.339 ;
        RECT 62.252 21.745 80 22.6 ;
        RECT 63.448 20.549 63.494 27.339 ;
        RECT 56.686 27.311 63.448 27.385 ;
        RECT 62.298 21.699 80 22.6 ;
        RECT 63.402 20.595 63.448 27.385 ;
        RECT 56.64 27.357 63.402 27.431 ;
        RECT 62.344 21.653 80 22.6 ;
        RECT 63.356 20.641 63.402 27.431 ;
        RECT 56.594 27.403 63.356 27.477 ;
        RECT 62.39 21.607 80 22.6 ;
        RECT 63.31 20.687 63.356 27.477 ;
        RECT 56.548 27.449 63.31 27.523 ;
        RECT 62.436 21.561 80 22.6 ;
        RECT 63.264 20.733 63.31 27.523 ;
        RECT 56.502 27.495 63.264 27.569 ;
        RECT 62.482 21.515 80 22.6 ;
        RECT 63.218 20.779 63.264 27.569 ;
        RECT 56.456 27.541 63.218 27.615 ;
        RECT 62.528 21.469 80 22.6 ;
        RECT 63.172 20.825 63.218 27.615 ;
        RECT 56.41 27.587 63.172 27.661 ;
        RECT 62.574 21.423 80 22.6 ;
        RECT 63.126 20.871 63.172 27.661 ;
        RECT 56.364 27.633 63.126 27.707 ;
        RECT 62.62 21.377 80 22.6 ;
        RECT 63.08 20.917 63.126 27.707 ;
        RECT 56.318 27.679 63.08 27.753 ;
        RECT 62.666 21.331 80 22.6 ;
        RECT 63.034 20.963 63.08 27.753 ;
        RECT 56.272 27.725 63.034 27.799 ;
        RECT 62.712 21.285 80 22.6 ;
        RECT 62.988 21.009 63.034 27.799 ;
        RECT 56.226 27.771 62.988 27.845 ;
        RECT 62.758 21.239 80 22.6 ;
        RECT 62.942 21.055 62.988 27.845 ;
        RECT 56.18 27.817 62.942 27.891 ;
        RECT 62.804 21.193 80 22.6 ;
        RECT 62.896 21.101 62.942 27.891 ;
        RECT 56.134 27.863 62.896 27.937 ;
        RECT 62.85 21.147 80 22.6 ;
        RECT 56.088 27.909 62.85 27.983 ;
        RECT 56.042 27.955 62.804 28.029 ;
        RECT 55.996 28.001 62.758 28.075 ;
        RECT 55.95 28.047 62.712 28.121 ;
        RECT 55.904 28.093 62.666 28.167 ;
        RECT 55.858 28.139 62.62 28.213 ;
        RECT 55.812 28.185 62.574 28.259 ;
        RECT 55.766 28.231 62.528 28.305 ;
        RECT 55.72 28.277 62.482 28.351 ;
        RECT 55.674 28.323 62.436 28.397 ;
        RECT 55.628 28.369 62.39 28.443 ;
        RECT 55.582 28.415 62.344 28.489 ;
        RECT 55.536 28.461 62.298 28.535 ;
        RECT 55.49 28.507 62.252 28.581 ;
        RECT 55.444 28.553 62.206 28.627 ;
        RECT 55.398 28.599 62.16 28.673 ;
        RECT 55.352 28.645 62.114 28.719 ;
        RECT 55.306 28.691 62.068 28.765 ;
        RECT 55.26 28.737 62.022 28.811 ;
        RECT 55.214 28.783 61.976 28.857 ;
        RECT 55.168 28.829 61.93 28.903 ;
        RECT 55.122 28.875 61.884 28.949 ;
        RECT 55.076 28.921 61.838 28.995 ;
        RECT 55.03 28.967 61.792 29.041 ;
        RECT 54.984 29.013 61.746 29.087 ;
        RECT 54.938 29.059 61.7 29.133 ;
        RECT 54.892 29.105 61.654 29.179 ;
        RECT 54.846 29.151 61.608 29.225 ;
        RECT 54.8 29.197 61.562 29.271 ;
        RECT 54.754 29.243 61.516 29.317 ;
        RECT 54.708 29.289 61.47 29.363 ;
        RECT 54.662 29.335 61.424 29.409 ;
        RECT 54.616 29.381 61.378 29.455 ;
        RECT 54.57 29.427 61.332 29.501 ;
        RECT 54.524 29.473 61.286 29.547 ;
        RECT 54.478 29.519 61.24 29.593 ;
        RECT 54.432 29.565 61.194 29.639 ;
        RECT 54.386 29.611 61.148 29.685 ;
        RECT 54.34 29.657 61.102 29.731 ;
        RECT 54.294 29.703 61.056 29.777 ;
        RECT 54.248 29.749 61.01 29.823 ;
        RECT 54.202 29.795 60.964 29.869 ;
        RECT 54.156 29.841 60.918 29.915 ;
        RECT 54.11 29.887 60.872 29.961 ;
        RECT 54.064 29.933 60.826 30.007 ;
        RECT 54.018 29.979 60.78 30.053 ;
        RECT 53.972 30.025 60.734 30.099 ;
        RECT 53.926 30.071 60.688 30.145 ;
        RECT 53.88 30.117 60.642 30.191 ;
        RECT 53.834 30.163 60.596 30.237 ;
        RECT 53.788 30.209 60.55 30.283 ;
        RECT 53.742 30.255 60.504 30.329 ;
        RECT 53.696 30.301 60.458 30.375 ;
        RECT 53.65 30.347 60.412 30.421 ;
        RECT 53.604 30.393 60.366 30.467 ;
        RECT 53.558 30.439 60.32 30.513 ;
        RECT 53.512 30.485 60.274 30.559 ;
        RECT 53.466 30.531 60.228 30.605 ;
        RECT 53.42 30.577 60.182 30.651 ;
        RECT 53.374 30.623 60.136 30.697 ;
        RECT 53.328 30.669 60.09 30.743 ;
        RECT 53.282 30.715 60.044 30.789 ;
        RECT 53.236 30.761 59.998 30.835 ;
        RECT 53.19 30.807 59.952 30.881 ;
        RECT 53.144 30.853 59.906 30.927 ;
        RECT 53.098 30.899 59.86 30.973 ;
        RECT 53.052 30.945 59.814 31.019 ;
        RECT 53.006 30.991 59.768 31.065 ;
        RECT 52.96 31.037 59.722 31.111 ;
        RECT 52.914 31.083 59.676 31.157 ;
        RECT 52.868 31.129 59.63 31.203 ;
        RECT 52.822 31.175 59.584 31.249 ;
        RECT 52.776 31.221 59.538 31.295 ;
        RECT 52.73 31.267 59.492 31.341 ;
        RECT 52.684 31.313 59.446 31.387 ;
        RECT 52.638 31.359 59.4 31.433 ;
        RECT 52.592 31.405 59.354 31.479 ;
        RECT 52.546 31.451 59.308 31.525 ;
        RECT 52.5 31.497 59.262 31.571 ;
        RECT 52.454 31.543 59.216 31.617 ;
        RECT 52.408 31.589 59.17 31.663 ;
        RECT 52.362 31.635 59.124 31.709 ;
        RECT 52.316 31.681 59.078 31.755 ;
        RECT 52.27 31.727 59.032 31.801 ;
        RECT 52.224 31.773 58.986 31.847 ;
        RECT 52.178 31.819 58.94 31.893 ;
        RECT 52.132 31.865 58.894 31.939 ;
        RECT 52.086 31.911 58.848 31.985 ;
        RECT 52.04 31.957 58.802 32.031 ;
        RECT 51.994 32.003 58.756 32.077 ;
        RECT 51.948 32.049 58.71 32.123 ;
        RECT 51.902 32.095 58.664 32.169 ;
        RECT 51.856 32.141 58.618 32.215 ;
        RECT 51.81 32.187 58.572 32.261 ;
        RECT 51.764 32.233 58.526 32.307 ;
        RECT 51.718 32.279 58.48 32.353 ;
        RECT 51.672 32.325 58.434 32.399 ;
        RECT 51.626 32.371 58.388 32.445 ;
        RECT 51.58 32.417 58.342 32.491 ;
        RECT 51.534 32.463 58.296 32.537 ;
        RECT 51.488 32.509 58.25 32.583 ;
        RECT 51.442 32.555 58.204 32.629 ;
        RECT 51.396 32.601 58.158 32.675 ;
        RECT 51.35 32.647 58.112 32.721 ;
        RECT 51.304 32.693 58.066 32.767 ;
        RECT 51.258 32.739 58.02 32.813 ;
        RECT 51.212 32.785 57.974 32.859 ;
        RECT 51.166 32.831 57.928 32.905 ;
        RECT 51.12 32.877 57.882 32.951 ;
        RECT 51.074 32.923 57.836 32.997 ;
        RECT 51.028 32.969 57.79 33.043 ;
        RECT 50.982 33.015 57.744 33.089 ;
        RECT 50.936 33.061 57.698 33.135 ;
        RECT 50.89 33.107 57.652 33.181 ;
        RECT 50.844 33.153 57.606 33.227 ;
        RECT 50.798 33.199 57.56 33.273 ;
        RECT 50.752 33.245 57.514 33.319 ;
        RECT 50.706 33.291 57.468 33.365 ;
        RECT 50.66 33.337 57.422 33.411 ;
        RECT 50.614 33.383 57.376 33.457 ;
        RECT 50.568 33.429 57.33 33.503 ;
        RECT 50.522 33.475 57.284 33.549 ;
        RECT 50.476 33.521 57.238 33.595 ;
        RECT 50.43 33.567 57.192 33.641 ;
        RECT 50.384 33.613 57.146 33.687 ;
        RECT 50.338 33.659 57.1 33.733 ;
        RECT 50.292 33.705 57.054 33.779 ;
        RECT 50.246 33.751 57.008 33.825 ;
        RECT 50.2 33.797 56.962 33.871 ;
        RECT 50.154 33.843 56.916 33.917 ;
        RECT 50.108 33.889 56.87 33.963 ;
        RECT 50.062 33.935 56.824 34.009 ;
        RECT 50.016 33.981 56.778 34.055 ;
        RECT 49.97 34.027 56.732 34.101 ;
        RECT 49.924 34.073 56.686 34.147 ;
        RECT 49.878 34.119 56.64 34.193 ;
        RECT 49.832 34.165 56.594 34.239 ;
        RECT 49.786 34.211 56.548 34.285 ;
        RECT 49.74 34.257 56.502 34.331 ;
        RECT 49.694 34.303 56.456 34.377 ;
        RECT 49.648 34.349 56.41 34.423 ;
        RECT 49.602 34.395 56.364 34.469 ;
        RECT 49.556 34.441 56.318 34.515 ;
        RECT 49.51 34.487 56.272 34.561 ;
        RECT 49.464 34.533 56.226 34.607 ;
        RECT 49.418 34.579 56.18 34.653 ;
        RECT 49.372 34.625 56.134 34.699 ;
        RECT 49.326 34.671 56.088 34.745 ;
        RECT 49.28 34.717 56.042 34.791 ;
        RECT 49.234 34.763 55.996 34.837 ;
        RECT 49.188 34.809 55.95 34.883 ;
        RECT 49.142 34.855 55.904 34.929 ;
        RECT 49.096 34.901 55.858 34.975 ;
        RECT 49.05 34.947 55.812 35.021 ;
        RECT 49.004 34.993 55.766 35.067 ;
        RECT 48.958 35.039 55.72 35.113 ;
        RECT 48.912 35.085 55.674 35.159 ;
        RECT 48.866 35.131 55.628 35.205 ;
        RECT 48.82 35.177 55.582 35.251 ;
        RECT 48.774 35.223 55.536 35.297 ;
        RECT 48.728 35.269 55.49 35.343 ;
        RECT 48.682 35.315 55.444 35.389 ;
        RECT 48.636 35.361 55.398 35.435 ;
        RECT 48.59 35.407 55.352 35.481 ;
        RECT 48.544 35.453 55.306 35.527 ;
        RECT 48.498 35.499 55.26 35.573 ;
        RECT 48.452 35.545 55.214 35.619 ;
        RECT 48.406 35.591 55.168 35.665 ;
        RECT 48.36 35.637 55.122 35.711 ;
        RECT 48.314 35.683 55.076 35.757 ;
        RECT 48.268 35.729 55.03 35.803 ;
        RECT 48.222 35.775 54.984 35.849 ;
        RECT 48.176 35.821 54.938 35.895 ;
        RECT 48.13 35.867 54.892 35.941 ;
        RECT 48.084 35.913 54.846 35.987 ;
        RECT 48.038 35.959 54.8 36.033 ;
        RECT 47.992 36.005 54.754 36.079 ;
        RECT 47.946 36.051 54.708 36.125 ;
        RECT 47.9 36.097 54.662 36.171 ;
        RECT 47.854 36.143 54.616 36.217 ;
        RECT 47.808 36.189 54.57 36.263 ;
        RECT 47.762 36.235 54.524 36.309 ;
        RECT 47.716 36.281 54.478 36.355 ;
        RECT 47.67 36.327 54.432 36.401 ;
        RECT 47.624 36.373 54.386 36.447 ;
        RECT 47.578 36.419 54.34 36.493 ;
        RECT 47.532 36.465 54.294 36.539 ;
        RECT 47.486 36.511 54.248 36.585 ;
        RECT 47.44 36.557 54.202 36.631 ;
        RECT 47.394 36.603 54.156 36.677 ;
        RECT 47.348 36.649 54.11 36.723 ;
        RECT 47.302 36.695 54.064 36.769 ;
        RECT 47.256 36.741 54.018 36.815 ;
        RECT 47.21 36.787 53.972 36.861 ;
        RECT 47.164 36.833 53.926 36.907 ;
        RECT 47.118 36.879 53.88 36.953 ;
        RECT 47.072 36.925 53.834 36.999 ;
        RECT 47.026 36.971 53.788 37.045 ;
        RECT 46.98 37.017 53.742 37.091 ;
        RECT 46.934 37.063 53.696 37.137 ;
        RECT 46.888 37.109 53.65 37.183 ;
        RECT 46.842 37.155 53.604 37.229 ;
        RECT 46.796 37.201 53.558 37.275 ;
        RECT 46.75 37.247 53.512 37.321 ;
        RECT 46.704 37.293 53.466 37.367 ;
        RECT 46.658 37.339 53.42 37.413 ;
        RECT 46.612 37.385 53.374 37.459 ;
        RECT 46.566 37.431 53.328 37.505 ;
        RECT 46.52 37.477 53.282 37.551 ;
        RECT 46.474 37.523 53.236 37.597 ;
        RECT 46.428 37.569 53.19 37.643 ;
        RECT 46.382 37.615 53.144 37.689 ;
        RECT 46.336 37.661 53.098 37.735 ;
        RECT 46.29 37.707 53.052 37.781 ;
        RECT 46.244 37.753 53.006 37.827 ;
        RECT 46.198 37.799 52.96 37.873 ;
        RECT 46.152 37.845 52.914 37.919 ;
        RECT 46.106 37.891 52.868 37.965 ;
        RECT 46.06 37.937 52.822 38.011 ;
        RECT 46.014 37.983 52.776 38.057 ;
        RECT 45.968 38.029 52.73 38.103 ;
        RECT 45.922 38.075 52.684 38.149 ;
        RECT 45.876 38.121 52.638 38.195 ;
        RECT 45.83 38.167 52.592 38.241 ;
        RECT 45.784 38.213 52.546 38.287 ;
        RECT 45.738 38.259 52.5 38.333 ;
        RECT 45.692 38.305 52.454 38.379 ;
        RECT 45.646 38.351 52.408 38.425 ;
        RECT 45.6 38.397 52.362 38.471 ;
        RECT 45.554 38.443 52.316 38.517 ;
        RECT 45.508 38.489 52.27 38.563 ;
        RECT 45.462 38.535 52.224 38.609 ;
        RECT 45.416 38.581 52.178 38.655 ;
        RECT 45.37 38.627 52.132 38.701 ;
        RECT 45.324 38.673 52.086 38.747 ;
        RECT 45.278 38.719 52.04 38.793 ;
        RECT 45.232 38.765 51.994 38.839 ;
        RECT 45.186 38.811 51.948 38.885 ;
        RECT 45.14 38.857 51.902 38.931 ;
        RECT 45.094 38.903 51.856 38.977 ;
        RECT 45.048 38.949 51.81 39.023 ;
        RECT 45.002 38.995 51.764 39.069 ;
        RECT 44.956 39.041 51.718 39.115 ;
        RECT 44.91 39.087 51.672 39.161 ;
        RECT 44.864 39.133 51.626 39.207 ;
        RECT 44.818 39.179 51.58 39.253 ;
        RECT 44.772 39.225 51.534 39.299 ;
        RECT 44.726 39.271 51.488 39.345 ;
        RECT 44.68 39.317 51.442 39.391 ;
        RECT 44.634 39.363 51.396 39.437 ;
        RECT 44.588 39.409 51.35 39.483 ;
        RECT 44.542 39.455 51.304 39.529 ;
        RECT 44.496 39.501 51.258 39.575 ;
        RECT 44.45 39.547 51.212 39.621 ;
        RECT 44.404 39.593 51.166 39.667 ;
        RECT 44.358 39.639 51.12 39.713 ;
        RECT 44.312 39.685 51.074 39.759 ;
        RECT 44.266 39.731 51.028 39.805 ;
        RECT 44.22 39.777 50.982 39.851 ;
        RECT 44.174 39.823 50.936 39.897 ;
        RECT 44.128 39.869 50.89 39.943 ;
        RECT 44.082 39.915 50.844 39.989 ;
        RECT 44.036 39.961 50.798 40.035 ;
        RECT 43.99 40.007 50.752 40.081 ;
        RECT 43.944 40.053 50.706 40.127 ;
        RECT 43.898 40.099 50.66 40.173 ;
        RECT 43.852 40.145 50.614 40.219 ;
        RECT 43.806 40.191 50.568 40.265 ;
        RECT 43.76 40.237 50.522 40.311 ;
        RECT 43.714 40.283 50.476 40.357 ;
        RECT 43.668 40.329 50.43 40.403 ;
        RECT 43.622 40.375 50.384 40.449 ;
        RECT 43.576 40.421 50.338 40.495 ;
        RECT 43.53 40.467 50.292 40.541 ;
        RECT 43.484 40.513 50.246 40.587 ;
        RECT 43.438 40.559 50.2 40.633 ;
        RECT 43.392 40.605 50.154 40.679 ;
        RECT 43.346 40.651 50.108 40.725 ;
        RECT 43.3 40.697 50.062 40.771 ;
        RECT 43.254 40.743 50.016 40.817 ;
        RECT 43.208 40.789 49.97 40.863 ;
        RECT 43.162 40.835 49.924 40.909 ;
        RECT 43.116 40.881 49.878 40.955 ;
        RECT 43.07 40.927 49.832 41.001 ;
        RECT 43.024 40.973 49.786 41.047 ;
        RECT 42.978 41.019 49.74 41.093 ;
        RECT 42.932 41.065 49.694 41.139 ;
        RECT 42.886 41.111 49.648 41.185 ;
        RECT 42.84 41.157 49.602 41.231 ;
        RECT 42.794 41.203 49.556 41.277 ;
        RECT 42.748 41.249 49.51 41.323 ;
        RECT 42.702 41.295 49.464 41.369 ;
        RECT 42.656 41.341 49.418 41.415 ;
        RECT 42.61 41.387 49.372 41.461 ;
        RECT 42.564 41.433 49.326 41.507 ;
        RECT 42.518 41.479 49.28 41.553 ;
        RECT 42.472 41.525 49.234 41.599 ;
        RECT 42.426 41.571 49.188 41.645 ;
        RECT 42.38 41.617 49.142 41.691 ;
        RECT 42.334 41.663 49.096 41.737 ;
        RECT 42.288 41.709 49.05 41.783 ;
        RECT 42.242 41.755 49.004 41.829 ;
        RECT 42.196 41.801 48.958 41.875 ;
        RECT 42.15 41.847 48.912 41.921 ;
        RECT 42.104 41.893 48.866 41.967 ;
        RECT 42.058 41.939 48.82 42.013 ;
        RECT 42.012 41.985 48.774 42.059 ;
        RECT 41.966 42.031 48.728 42.105 ;
        RECT 41.92 42.077 48.682 42.151 ;
        RECT 41.874 42.123 48.636 42.197 ;
        RECT 41.828 42.169 48.59 42.243 ;
        RECT 41.782 42.215 48.544 42.289 ;
        RECT 41.736 42.261 48.498 42.335 ;
        RECT 41.69 42.307 48.452 42.381 ;
        RECT 41.644 42.353 48.406 42.427 ;
        RECT 41.598 42.399 48.36 42.473 ;
        RECT 41.552 42.445 48.314 42.519 ;
        RECT 41.506 42.491 48.268 42.565 ;
        RECT 41.46 42.537 48.222 42.611 ;
        RECT 41.414 42.583 48.176 42.657 ;
        RECT 41.368 42.629 48.13 42.703 ;
        RECT 41.322 42.675 48.084 42.749 ;
        RECT 41.276 42.721 48.038 42.795 ;
        RECT 41.23 42.767 47.992 42.841 ;
        RECT 41.184 42.813 47.946 42.887 ;
        RECT 41.138 42.859 47.9 42.933 ;
        RECT 41.092 42.905 47.854 42.979 ;
        RECT 41.046 42.951 47.808 43.025 ;
        RECT 41 42.997 47.762 43.071 ;
        RECT 40.954 43.043 47.716 43.117 ;
        RECT 40.908 43.089 47.67 43.163 ;
        RECT 40.862 43.135 47.624 43.209 ;
        RECT 40.816 43.181 47.578 43.255 ;
        RECT 40.77 43.227 47.532 43.301 ;
        RECT 40.724 43.273 47.486 43.347 ;
        RECT 40.678 43.319 47.44 43.393 ;
        RECT 40.632 43.365 47.394 43.439 ;
        RECT 40.586 43.411 47.348 43.485 ;
        RECT 40.54 43.457 47.302 43.531 ;
        RECT 40.494 43.503 47.256 43.577 ;
        RECT 40.448 43.549 47.21 43.623 ;
        RECT 40.402 43.595 47.164 43.669 ;
        RECT 40.356 43.641 47.118 43.715 ;
        RECT 40.31 43.687 47.072 43.761 ;
        RECT 40.264 43.733 47.026 43.807 ;
        RECT 40.218 43.779 46.98 43.853 ;
        RECT 40.172 43.825 46.934 43.899 ;
        RECT 40.126 43.871 46.888 43.945 ;
        RECT 40.08 43.917 46.842 43.991 ;
        RECT 40.034 43.963 46.796 44.037 ;
        RECT 39.988 44.009 46.75 44.083 ;
        RECT 39.942 44.055 46.704 44.129 ;
        RECT 39.896 44.101 46.658 44.175 ;
        RECT 39.85 44.147 46.612 44.221 ;
        RECT 39.804 44.193 46.566 44.267 ;
        RECT 39.758 44.239 46.52 44.313 ;
        RECT 39.712 44.285 46.474 44.359 ;
        RECT 39.666 44.331 46.428 44.405 ;
        RECT 39.62 44.377 46.382 44.451 ;
        RECT 39.574 44.423 46.336 44.497 ;
        RECT 39.528 44.469 46.29 44.543 ;
        RECT 39.482 44.515 46.244 44.589 ;
        RECT 39.436 44.561 46.198 44.635 ;
        RECT 39.39 44.607 46.152 44.681 ;
        RECT 39.344 44.653 46.106 44.727 ;
        RECT 39.298 44.699 46.06 44.773 ;
        RECT 39.252 44.745 46.014 44.819 ;
        RECT 39.206 44.791 45.968 44.865 ;
        RECT 39.16 44.837 45.922 44.911 ;
        RECT 39.114 44.883 45.876 44.957 ;
        RECT 39.068 44.929 45.83 45.003 ;
        RECT 39.022 44.975 45.784 45.049 ;
        RECT 38.976 45.021 45.738 45.095 ;
        RECT 38.93 45.067 45.692 45.141 ;
        RECT 38.884 45.113 45.646 45.187 ;
        RECT 38.838 45.159 45.6 45.233 ;
        RECT 38.792 45.205 45.554 45.279 ;
        RECT 38.746 45.251 45.508 45.325 ;
        RECT 38.7 45.297 45.462 45.371 ;
        RECT 38.654 45.343 45.416 45.417 ;
        RECT 38.608 45.389 45.37 45.463 ;
        RECT 38.562 45.435 45.324 45.509 ;
        RECT 38.516 45.481 45.278 45.555 ;
        RECT 38.47 45.527 45.232 45.601 ;
        RECT 38.424 45.573 45.186 45.647 ;
        RECT 38.378 45.619 45.14 45.693 ;
        RECT 38.332 45.665 45.094 45.739 ;
        RECT 38.286 45.711 45.048 45.785 ;
        RECT 38.24 45.757 45.002 45.831 ;
        RECT 38.194 45.803 44.956 45.877 ;
        RECT 38.148 45.849 44.91 45.923 ;
        RECT 38.102 45.895 44.864 45.969 ;
        RECT 38.056 45.941 44.818 46.015 ;
        RECT 38.01 45.987 44.772 46.061 ;
        RECT 37.964 46.033 44.726 46.107 ;
        RECT 37.918 46.079 44.68 46.153 ;
        RECT 37.872 46.125 44.634 46.199 ;
        RECT 37.826 46.171 44.588 46.245 ;
        RECT 37.78 46.217 44.542 46.291 ;
        RECT 37.734 46.263 44.496 46.337 ;
        RECT 37.688 46.309 44.45 46.383 ;
        RECT 37.642 46.355 44.404 46.429 ;
        RECT 37.596 46.401 44.358 46.475 ;
        RECT 37.55 46.447 44.312 46.521 ;
        RECT 37.504 46.493 44.266 46.567 ;
        RECT 37.458 46.539 44.22 46.613 ;
        RECT 37.412 46.585 44.174 46.659 ;
        RECT 37.366 46.631 44.128 46.705 ;
        RECT 37.32 46.677 44.082 46.751 ;
        RECT 37.274 46.723 44.036 46.797 ;
        RECT 37.228 46.769 43.99 46.843 ;
        RECT 37.182 46.815 43.944 46.889 ;
        RECT 37.136 46.861 43.898 46.935 ;
        RECT 37.09 46.907 43.852 46.981 ;
        RECT 37.044 46.953 43.806 47.027 ;
        RECT 36.998 46.999 43.76 47.073 ;
        RECT 36.952 47.045 43.714 47.119 ;
        RECT 36.906 47.091 43.668 47.165 ;
        RECT 36.86 47.137 43.622 47.211 ;
        RECT 36.814 47.183 43.576 47.257 ;
        RECT 36.768 47.229 43.53 47.303 ;
        RECT 36.722 47.275 43.484 47.349 ;
        RECT 36.676 47.321 43.438 47.395 ;
        RECT 36.63 47.367 43.392 47.441 ;
        RECT 36.584 47.413 43.346 47.487 ;
        RECT 36.538 47.459 43.3 47.533 ;
        RECT 36.492 47.505 43.254 47.579 ;
        RECT 36.446 47.551 43.208 47.625 ;
        RECT 36.4 47.597 43.162 47.671 ;
        RECT 36.354 47.643 43.116 47.717 ;
        RECT 36.308 47.689 43.07 47.763 ;
        RECT 36.262 47.735 43.024 47.809 ;
        RECT 36.216 47.781 42.978 47.855 ;
        RECT 36.17 47.827 42.932 47.901 ;
        RECT 36.124 47.873 42.886 47.947 ;
        RECT 36.078 47.919 42.84 47.993 ;
        RECT 36.032 47.965 42.794 48.039 ;
        RECT 35.986 48.011 42.748 48.085 ;
        RECT 35.94 48.057 42.702 48.131 ;
        RECT 35.894 48.103 42.656 48.177 ;
        RECT 35.848 48.149 42.61 48.223 ;
        RECT 35.802 48.195 42.564 48.269 ;
        RECT 35.756 48.241 42.518 48.315 ;
        RECT 35.71 48.287 42.472 48.361 ;
        RECT 35.664 48.333 42.426 48.407 ;
        RECT 35.618 48.379 42.38 48.453 ;
        RECT 35.572 48.425 42.334 48.499 ;
        RECT 35.526 48.471 42.288 48.545 ;
        RECT 35.48 48.517 42.242 48.591 ;
        RECT 35.434 48.563 42.196 48.637 ;
        RECT 35.388 48.609 42.15 48.683 ;
        RECT 35.342 48.655 42.104 48.729 ;
        RECT 35.296 48.701 42.058 48.775 ;
        RECT 35.25 48.747 42.012 48.821 ;
        RECT 35.204 48.793 41.966 48.867 ;
        RECT 35.158 48.839 41.92 48.913 ;
        RECT 35.112 48.885 41.874 48.959 ;
        RECT 35.066 48.931 41.828 49.005 ;
        RECT 35.02 48.977 41.782 49.051 ;
        RECT 34.974 49.023 41.736 49.097 ;
        RECT 34.928 49.069 41.69 49.143 ;
        RECT 34.882 49.115 41.644 49.189 ;
        RECT 34.836 49.161 41.598 49.235 ;
        RECT 34.79 49.207 41.552 49.281 ;
        RECT 34.744 49.253 41.506 49.327 ;
        RECT 34.698 49.299 41.46 49.373 ;
        RECT 34.652 49.345 41.414 49.419 ;
        RECT 34.606 49.391 41.368 49.465 ;
        RECT 34.56 49.437 41.322 49.511 ;
        RECT 34.514 49.483 41.276 49.557 ;
        RECT 34.468 49.529 41.23 49.603 ;
        RECT 34.422 49.575 41.184 49.649 ;
        RECT 34.376 49.621 41.138 49.695 ;
        RECT 34.33 49.667 41.092 49.741 ;
        RECT 34.284 49.713 41.046 49.787 ;
        RECT 34.238 49.759 41 49.833 ;
        RECT 34.192 49.805 40.954 49.879 ;
        RECT 34.146 49.851 40.908 49.925 ;
        RECT 34.1 49.897 40.862 49.971 ;
        RECT 34.054 49.943 40.816 50.017 ;
        RECT 34.008 49.989 40.77 50.063 ;
        RECT 33.962 50.035 40.724 50.109 ;
        RECT 33.916 50.081 40.678 50.155 ;
        RECT 33.87 50.127 40.632 50.201 ;
        RECT 33.824 50.173 40.586 50.247 ;
        RECT 33.778 50.219 40.54 50.293 ;
        RECT 33.732 50.265 40.494 50.339 ;
        RECT 33.686 50.311 40.448 50.385 ;
        RECT 33.64 50.357 40.402 50.431 ;
        RECT 33.594 50.403 40.356 50.477 ;
        RECT 33.548 50.449 40.31 50.523 ;
        RECT 33.502 50.495 40.264 50.569 ;
        RECT 33.456 50.541 40.218 50.615 ;
        RECT 33.41 50.587 40.172 50.661 ;
        RECT 33.364 50.633 40.126 50.707 ;
        RECT 33.318 50.679 40.08 50.753 ;
        RECT 33.272 50.725 40.034 50.799 ;
        RECT 33.226 50.771 39.988 50.845 ;
        RECT 33.18 50.817 39.942 50.891 ;
        RECT 33.134 50.863 39.896 50.937 ;
        RECT 33.088 50.909 39.85 50.983 ;
        RECT 33.042 50.955 39.804 51.029 ;
        RECT 32.996 51.001 39.758 51.075 ;
        RECT 32.95 51.047 39.712 51.121 ;
        RECT 32.904 51.093 39.666 51.167 ;
        RECT 32.858 51.139 39.62 51.213 ;
        RECT 32.812 51.185 39.574 51.259 ;
        RECT 32.766 51.231 39.528 51.305 ;
        RECT 32.72 51.277 39.482 51.351 ;
        RECT 32.674 51.323 39.436 51.397 ;
        RECT 32.628 51.369 39.39 51.443 ;
        RECT 32.582 51.415 39.344 51.489 ;
        RECT 32.536 51.461 39.298 51.535 ;
        RECT 32.49 51.507 39.252 51.581 ;
        RECT 32.444 51.553 39.206 51.627 ;
        RECT 32.398 51.599 39.16 51.673 ;
        RECT 32.352 51.645 39.114 51.719 ;
        RECT 32.306 51.691 39.068 51.765 ;
        RECT 32.26 51.737 39.022 51.811 ;
        RECT 32.214 51.783 38.976 51.857 ;
        RECT 32.168 51.829 38.93 51.903 ;
        RECT 32.122 51.875 38.884 51.949 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 78.01 67.4 80 72.206 ;
        RECT 71.264 74.123 78.01 74.197 ;
        RECT 71.31 74.077 78.056 74.167 ;
        RECT 77.996 67.407 78.01 74.197 ;
        RECT 71.218 74.169 77.996 74.227 ;
        RECT 71.356 74.031 78.102 74.121 ;
        RECT 77.95 67.437 77.996 74.227 ;
        RECT 71.172 74.215 77.95 74.273 ;
        RECT 71.402 73.985 78.148 74.075 ;
        RECT 77.904 67.483 77.95 74.273 ;
        RECT 71.126 74.261 77.904 74.319 ;
        RECT 71.448 73.939 78.194 74.029 ;
        RECT 77.858 67.529 77.904 74.319 ;
        RECT 71.08 74.307 77.858 74.365 ;
        RECT 71.494 73.893 78.24 73.983 ;
        RECT 77.812 67.575 77.858 74.365 ;
        RECT 71.034 74.353 77.812 74.411 ;
        RECT 71.54 73.847 78.286 73.937 ;
        RECT 77.766 67.621 77.812 74.411 ;
        RECT 70.988 74.399 77.766 74.457 ;
        RECT 71.586 73.801 78.332 73.891 ;
        RECT 77.72 67.667 77.766 74.457 ;
        RECT 70.942 74.445 77.72 74.503 ;
        RECT 71.632 73.755 78.378 73.845 ;
        RECT 77.674 67.713 77.72 74.503 ;
        RECT 70.896 74.491 77.674 74.549 ;
        RECT 71.678 73.709 78.424 73.799 ;
        RECT 77.628 67.759 77.674 74.549 ;
        RECT 70.85 74.537 77.628 74.595 ;
        RECT 71.724 73.663 78.47 73.753 ;
        RECT 77.582 67.805 77.628 74.595 ;
        RECT 70.804 74.583 77.582 74.641 ;
        RECT 71.77 73.617 78.516 73.707 ;
        RECT 77.536 67.851 77.582 74.641 ;
        RECT 70.758 74.629 77.536 74.687 ;
        RECT 71.816 73.571 78.562 73.661 ;
        RECT 77.49 67.897 77.536 74.687 ;
        RECT 70.712 74.675 77.49 74.733 ;
        RECT 71.862 73.525 78.608 73.615 ;
        RECT 77.444 67.943 77.49 74.733 ;
        RECT 70.666 74.721 77.444 74.779 ;
        RECT 71.908 73.479 78.654 73.569 ;
        RECT 77.398 67.989 77.444 74.779 ;
        RECT 70.62 74.767 77.398 74.825 ;
        RECT 71.954 73.433 78.7 73.523 ;
        RECT 77.352 68.035 77.398 74.825 ;
        RECT 70.574 74.813 77.352 74.871 ;
        RECT 72 73.387 78.746 73.477 ;
        RECT 77.306 68.081 77.352 74.871 ;
        RECT 70.528 74.859 77.306 74.917 ;
        RECT 72.046 73.341 78.792 73.431 ;
        RECT 77.26 68.127 77.306 74.917 ;
        RECT 70.482 74.905 77.26 74.963 ;
        RECT 72.092 73.295 78.838 73.385 ;
        RECT 77.214 68.173 77.26 74.963 ;
        RECT 70.436 74.951 77.214 75.009 ;
        RECT 72.138 73.249 78.884 73.339 ;
        RECT 77.168 68.219 77.214 75.009 ;
        RECT 70.39 74.997 77.168 75.055 ;
        RECT 72.184 73.218 78.93 73.293 ;
        RECT 77.122 68.265 77.168 75.055 ;
        RECT 70.344 75.043 77.122 75.101 ;
        RECT 72.2 73.187 78.976 73.247 ;
        RECT 77.076 68.311 77.122 75.101 ;
        RECT 70.298 75.089 77.076 75.147 ;
        RECT 72.246 73.141 79.022 73.201 ;
        RECT 77.03 68.357 77.076 75.147 ;
        RECT 70.252 75.135 77.03 75.193 ;
        RECT 72.292 73.095 79.068 73.155 ;
        RECT 76.984 68.403 77.03 75.193 ;
        RECT 70.206 75.181 76.984 75.239 ;
        RECT 72.338 73.049 79.114 73.109 ;
        RECT 76.938 68.449 76.984 75.239 ;
        RECT 70.16 75.227 76.938 75.285 ;
        RECT 72.384 73.003 79.16 73.063 ;
        RECT 76.892 68.495 76.938 75.285 ;
        RECT 70.114 75.273 76.892 75.331 ;
        RECT 72.43 72.957 79.206 73.017 ;
        RECT 76.846 68.541 76.892 75.331 ;
        RECT 70.068 75.319 76.846 75.377 ;
        RECT 72.476 72.911 79.252 72.971 ;
        RECT 76.8 68.587 76.846 75.377 ;
        RECT 70.022 75.365 76.8 75.423 ;
        RECT 72.522 72.865 79.298 72.925 ;
        RECT 76.754 68.633 76.8 75.423 ;
        RECT 69.976 75.411 76.754 75.469 ;
        RECT 72.568 72.819 79.344 72.879 ;
        RECT 76.708 68.679 76.754 75.469 ;
        RECT 69.93 75.457 76.708 75.515 ;
        RECT 72.614 72.773 79.39 72.833 ;
        RECT 76.662 68.725 76.708 75.515 ;
        RECT 69.884 75.503 76.662 75.561 ;
        RECT 72.66 72.727 79.436 72.787 ;
        RECT 76.616 68.771 76.662 75.561 ;
        RECT 69.838 75.549 76.616 75.607 ;
        RECT 72.706 72.681 79.482 72.741 ;
        RECT 76.57 68.817 76.616 75.607 ;
        RECT 69.792 75.595 76.57 75.653 ;
        RECT 72.752 72.635 79.528 72.695 ;
        RECT 76.524 68.863 76.57 75.653 ;
        RECT 69.746 75.641 76.524 75.699 ;
        RECT 72.798 72.589 79.574 72.649 ;
        RECT 76.478 68.909 76.524 75.699 ;
        RECT 69.7 75.687 76.478 75.745 ;
        RECT 72.844 72.543 79.62 72.603 ;
        RECT 76.432 68.955 76.478 75.745 ;
        RECT 69.654 75.733 76.432 75.791 ;
        RECT 72.89 72.497 79.666 72.557 ;
        RECT 76.386 69.001 76.432 75.791 ;
        RECT 69.608 75.779 76.386 75.837 ;
        RECT 72.936 72.451 79.712 72.511 ;
        RECT 76.34 69.047 76.386 75.837 ;
        RECT 69.562 75.825 76.34 75.883 ;
        RECT 72.982 72.405 79.758 72.465 ;
        RECT 76.294 69.093 76.34 75.883 ;
        RECT 69.516 75.871 76.294 75.929 ;
        RECT 73.028 72.359 79.804 72.419 ;
        RECT 76.248 69.139 76.294 75.929 ;
        RECT 69.47 75.917 76.248 75.975 ;
        RECT 73.074 72.313 79.85 72.373 ;
        RECT 76.202 69.185 76.248 75.975 ;
        RECT 69.424 75.963 76.202 76.021 ;
        RECT 73.12 72.267 79.896 72.327 ;
        RECT 76.156 69.231 76.202 76.021 ;
        RECT 69.378 76.009 76.156 76.067 ;
        RECT 73.166 72.221 79.942 72.281 ;
        RECT 76.11 69.277 76.156 76.067 ;
        RECT 69.332 76.055 76.11 76.113 ;
        RECT 73.212 72.175 79.988 72.235 ;
        RECT 76.064 69.323 76.11 76.113 ;
        RECT 69.286 76.101 76.064 76.159 ;
        RECT 73.258 72.129 80 72.206 ;
        RECT 76.018 69.369 76.064 76.159 ;
        RECT 69.24 76.147 76.018 76.205 ;
        RECT 73.304 72.083 80 72.206 ;
        RECT 75.972 69.415 76.018 76.205 ;
        RECT 69.194 76.193 75.972 76.251 ;
        RECT 73.35 72.037 80 72.206 ;
        RECT 75.926 69.461 75.972 76.251 ;
        RECT 69.148 76.239 75.926 76.297 ;
        RECT 73.396 71.991 80 72.206 ;
        RECT 75.88 69.507 75.926 76.297 ;
        RECT 69.102 76.285 75.88 76.343 ;
        RECT 73.442 71.945 80 72.206 ;
        RECT 75.834 69.553 75.88 76.343 ;
        RECT 69.056 76.331 75.834 76.389 ;
        RECT 73.488 71.899 80 72.206 ;
        RECT 75.788 69.599 75.834 76.389 ;
        RECT 69.01 76.377 75.788 76.435 ;
        RECT 73.534 71.853 80 72.206 ;
        RECT 75.742 69.645 75.788 76.435 ;
        RECT 68.964 76.423 75.742 76.481 ;
        RECT 73.58 71.807 80 72.206 ;
        RECT 75.696 69.691 75.742 76.481 ;
        RECT 68.918 76.469 75.696 76.527 ;
        RECT 73.626 71.761 80 72.206 ;
        RECT 75.65 69.737 75.696 76.527 ;
        RECT 68.872 76.515 75.65 76.573 ;
        RECT 73.672 71.715 80 72.206 ;
        RECT 75.604 69.783 75.65 76.573 ;
        RECT 68.826 76.561 75.604 76.619 ;
        RECT 73.718 71.669 80 72.206 ;
        RECT 75.558 69.829 75.604 76.619 ;
        RECT 68.78 76.607 75.558 76.665 ;
        RECT 73.764 71.623 80 72.206 ;
        RECT 75.512 69.875 75.558 76.665 ;
        RECT 68.734 76.653 75.512 76.711 ;
        RECT 73.81 71.577 80 72.206 ;
        RECT 75.466 69.921 75.512 76.711 ;
        RECT 68.688 76.699 75.466 76.757 ;
        RECT 73.856 71.531 80 72.206 ;
        RECT 75.42 69.967 75.466 76.757 ;
        RECT 68.642 76.745 75.42 76.803 ;
        RECT 73.902 71.485 80 72.206 ;
        RECT 75.374 70.013 75.42 76.803 ;
        RECT 68.596 76.791 75.374 76.849 ;
        RECT 73.948 71.439 80 72.206 ;
        RECT 75.328 70.059 75.374 76.849 ;
        RECT 68.55 76.837 75.328 76.895 ;
        RECT 73.994 71.393 80 72.206 ;
        RECT 75.282 70.105 75.328 76.895 ;
        RECT 68.504 76.883 75.282 76.941 ;
        RECT 74.04 71.347 80 72.206 ;
        RECT 75.236 70.151 75.282 76.941 ;
        RECT 68.458 76.929 75.236 76.987 ;
        RECT 74.086 71.301 80 72.206 ;
        RECT 75.19 70.197 75.236 76.987 ;
        RECT 68.412 76.975 75.19 77.033 ;
        RECT 74.132 71.255 80 72.206 ;
        RECT 75.144 70.243 75.19 77.033 ;
        RECT 68.366 77.021 75.144 77.079 ;
        RECT 74.178 71.209 80 72.206 ;
        RECT 75.098 70.289 75.144 77.079 ;
        RECT 68.32 77.067 75.098 77.125 ;
        RECT 74.224 71.163 80 72.206 ;
        RECT 75.052 70.335 75.098 77.125 ;
        RECT 68.274 77.113 75.052 77.171 ;
        RECT 74.27 71.117 80 72.206 ;
        RECT 75.006 70.381 75.052 77.171 ;
        RECT 68.228 77.159 75.006 77.217 ;
        RECT 74.316 71.071 80 72.206 ;
        RECT 74.96 70.427 75.006 77.217 ;
        RECT 68.182 77.205 74.96 77.263 ;
        RECT 74.362 71.025 80 72.206 ;
        RECT 74.914 70.473 74.96 77.263 ;
        RECT 68.136 77.251 74.914 77.309 ;
        RECT 74.408 70.979 80 72.206 ;
        RECT 74.868 70.519 74.914 77.309 ;
        RECT 68.09 77.297 74.868 77.355 ;
        RECT 74.454 70.933 80 72.206 ;
        RECT 74.822 70.565 74.868 77.355 ;
        RECT 68.044 77.343 74.822 77.401 ;
        RECT 74.5 70.887 80 72.206 ;
        RECT 74.776 70.611 74.822 77.401 ;
        RECT 67.998 77.389 74.776 77.447 ;
        RECT 74.546 70.841 80 72.206 ;
        RECT 74.73 70.657 74.776 77.447 ;
        RECT 67.952 77.435 74.73 77.493 ;
        RECT 74.592 70.795 80 72.206 ;
        RECT 74.684 70.703 74.73 77.493 ;
        RECT 67.906 77.481 74.684 77.539 ;
        RECT 74.638 70.749 80 72.206 ;
        RECT 67.86 77.527 74.638 77.585 ;
        RECT 67.814 77.573 74.592 77.631 ;
        RECT 67.768 77.619 74.546 77.677 ;
        RECT 67.722 77.665 74.5 77.723 ;
        RECT 67.676 77.711 74.454 77.769 ;
        RECT 67.63 77.757 74.408 77.815 ;
        RECT 67.584 77.803 74.362 77.861 ;
        RECT 67.538 77.849 74.316 77.907 ;
        RECT 67.492 77.895 74.27 77.953 ;
        RECT 67.446 77.941 74.224 77.999 ;
        RECT 67.4 77.987 74.178 78.045 ;
        RECT 67.4 77.987 74.132 78.091 ;
        RECT 67.4 77.987 74.086 78.137 ;
        RECT 67.4 77.987 74.04 78.183 ;
        RECT 67.4 77.987 73.994 78.229 ;
        RECT 67.4 77.987 73.948 78.275 ;
        RECT 67.4 77.987 73.902 78.321 ;
        RECT 67.4 77.987 73.856 78.367 ;
        RECT 67.4 77.987 73.81 78.413 ;
        RECT 67.4 77.987 73.764 78.459 ;
        RECT 67.4 77.987 73.718 78.505 ;
        RECT 67.4 77.987 73.672 78.551 ;
        RECT 67.4 77.987 73.626 78.597 ;
        RECT 67.4 77.987 73.58 78.643 ;
        RECT 67.4 77.987 73.534 78.689 ;
        RECT 67.4 77.987 73.488 78.735 ;
        RECT 67.4 77.987 73.442 78.781 ;
        RECT 67.4 77.987 73.396 78.827 ;
        RECT 67.4 77.987 73.35 78.873 ;
        RECT 67.4 77.987 73.304 78.919 ;
        RECT 67.4 77.987 73.258 78.965 ;
        RECT 67.4 77.987 73.212 79.011 ;
        RECT 67.4 77.987 73.166 79.057 ;
        RECT 67.4 77.987 73.12 79.103 ;
        RECT 67.4 77.987 73.074 79.149 ;
        RECT 67.4 77.987 73.028 79.195 ;
        RECT 67.4 77.987 72.982 79.241 ;
        RECT 67.4 77.987 72.936 79.287 ;
        RECT 67.4 77.987 72.89 79.333 ;
        RECT 67.4 77.987 72.844 79.379 ;
        RECT 67.4 77.987 72.798 79.425 ;
        RECT 67.4 77.987 72.752 79.471 ;
        RECT 67.4 77.987 72.706 79.517 ;
        RECT 67.4 77.987 72.66 79.563 ;
        RECT 67.4 77.987 72.614 79.609 ;
        RECT 67.4 77.987 72.568 79.655 ;
        RECT 67.4 77.987 72.522 79.701 ;
        RECT 67.4 77.987 72.476 79.747 ;
        RECT 67.4 77.987 72.43 79.793 ;
        RECT 67.4 77.987 72.384 79.839 ;
        RECT 67.4 77.987 72.338 79.885 ;
        RECT 67.4 77.987 72.292 79.931 ;
        RECT 67.4 77.987 72.246 79.977 ;
        RECT 67.4 77.987 72.2 80 ;
    END
    PORT
      LAYER QB ;
        RECT 70.3 48.8 80 53.6 ;
        RECT 65.514 53.563 72.29 53.606 ;
        RECT 63.536 55.541 70.3 55.591 ;
        RECT 63.582 55.495 70.346 55.567 ;
        RECT 70.298 48.801 70.3 55.591 ;
        RECT 63.628 55.449 70.392 55.521 ;
        RECT 70.252 48.825 70.298 55.615 ;
        RECT 63.49 55.587 70.252 55.661 ;
        RECT 63.674 55.403 70.438 55.475 ;
        RECT 70.206 48.871 70.252 55.661 ;
        RECT 63.444 55.633 70.206 55.707 ;
        RECT 63.72 55.357 70.484 55.429 ;
        RECT 70.16 48.917 70.206 55.707 ;
        RECT 63.398 55.679 70.16 55.753 ;
        RECT 63.766 55.311 70.53 55.383 ;
        RECT 70.114 48.963 70.16 55.753 ;
        RECT 63.352 55.725 70.114 55.799 ;
        RECT 63.812 55.265 70.576 55.337 ;
        RECT 70.068 49.009 70.114 55.799 ;
        RECT 63.306 55.771 70.068 55.845 ;
        RECT 63.858 55.219 70.622 55.291 ;
        RECT 70.022 49.055 70.068 55.845 ;
        RECT 63.26 55.817 70.022 55.891 ;
        RECT 63.904 55.173 70.668 55.245 ;
        RECT 69.976 49.101 70.022 55.891 ;
        RECT 63.214 55.863 69.976 55.937 ;
        RECT 63.95 55.127 70.714 55.199 ;
        RECT 69.93 49.147 69.976 55.937 ;
        RECT 63.168 55.909 69.93 55.983 ;
        RECT 63.996 55.081 70.76 55.153 ;
        RECT 69.884 49.193 69.93 55.983 ;
        RECT 63.122 55.955 69.884 56.029 ;
        RECT 64.042 55.035 70.806 55.107 ;
        RECT 69.838 49.239 69.884 56.029 ;
        RECT 63.076 56.001 69.838 56.075 ;
        RECT 64.088 54.989 70.852 55.061 ;
        RECT 69.792 49.285 69.838 56.075 ;
        RECT 63.03 56.047 69.792 56.121 ;
        RECT 64.134 54.943 70.898 55.015 ;
        RECT 69.746 49.331 69.792 56.121 ;
        RECT 62.984 56.093 69.746 56.167 ;
        RECT 64.18 54.897 70.944 54.969 ;
        RECT 69.7 49.377 69.746 56.167 ;
        RECT 62.938 56.139 69.7 56.213 ;
        RECT 64.226 54.851 70.99 54.923 ;
        RECT 69.654 49.423 69.7 56.213 ;
        RECT 62.892 56.185 69.654 56.259 ;
        RECT 64.272 54.805 71.036 54.877 ;
        RECT 69.608 49.469 69.654 56.259 ;
        RECT 62.846 56.231 69.608 56.305 ;
        RECT 64.318 54.759 71.082 54.831 ;
        RECT 69.562 49.515 69.608 56.305 ;
        RECT 62.8 56.277 69.562 56.351 ;
        RECT 64.364 54.713 71.128 54.785 ;
        RECT 69.516 49.561 69.562 56.351 ;
        RECT 62.754 56.323 69.516 56.397 ;
        RECT 64.41 54.667 71.174 54.739 ;
        RECT 69.47 49.607 69.516 56.397 ;
        RECT 62.708 56.369 69.47 56.443 ;
        RECT 64.456 54.621 71.22 54.693 ;
        RECT 69.424 49.653 69.47 56.443 ;
        RECT 62.662 56.415 69.424 56.489 ;
        RECT 64.502 54.575 71.266 54.647 ;
        RECT 69.378 49.699 69.424 56.489 ;
        RECT 62.616 56.461 69.378 56.535 ;
        RECT 64.548 54.529 71.312 54.601 ;
        RECT 69.332 49.745 69.378 56.535 ;
        RECT 62.57 56.507 69.332 56.581 ;
        RECT 64.594 54.483 71.358 54.555 ;
        RECT 69.286 49.791 69.332 56.581 ;
        RECT 62.524 56.553 69.286 56.627 ;
        RECT 64.64 54.437 71.404 54.509 ;
        RECT 69.24 49.837 69.286 56.627 ;
        RECT 62.478 56.599 69.24 56.673 ;
        RECT 64.686 54.391 71.45 54.463 ;
        RECT 69.194 49.883 69.24 56.673 ;
        RECT 62.432 56.645 69.194 56.719 ;
        RECT 64.732 54.345 71.496 54.417 ;
        RECT 69.148 49.929 69.194 56.719 ;
        RECT 62.386 56.691 69.148 56.765 ;
        RECT 64.778 54.299 71.542 54.371 ;
        RECT 69.102 49.975 69.148 56.765 ;
        RECT 62.34 56.737 69.102 56.811 ;
        RECT 64.824 54.253 71.588 54.325 ;
        RECT 69.056 50.021 69.102 56.811 ;
        RECT 62.294 56.783 69.056 56.857 ;
        RECT 64.87 54.207 71.634 54.279 ;
        RECT 69.01 50.067 69.056 56.857 ;
        RECT 62.248 56.829 69.01 56.903 ;
        RECT 64.916 54.161 71.68 54.233 ;
        RECT 68.964 50.113 69.01 56.903 ;
        RECT 62.202 56.875 68.964 56.949 ;
        RECT 64.962 54.115 71.726 54.187 ;
        RECT 68.918 50.159 68.964 56.949 ;
        RECT 62.156 56.921 68.918 56.995 ;
        RECT 65.008 54.069 71.772 54.141 ;
        RECT 68.872 50.205 68.918 56.995 ;
        RECT 62.11 56.967 68.872 57.041 ;
        RECT 65.054 54.023 71.818 54.095 ;
        RECT 68.826 50.251 68.872 57.041 ;
        RECT 62.064 57.013 68.826 57.087 ;
        RECT 65.1 53.977 71.864 54.049 ;
        RECT 68.78 50.297 68.826 57.087 ;
        RECT 62.018 57.059 68.78 57.133 ;
        RECT 65.146 53.931 71.91 54.003 ;
        RECT 68.734 50.343 68.78 57.133 ;
        RECT 61.972 57.105 68.734 57.179 ;
        RECT 65.192 53.885 71.956 53.957 ;
        RECT 68.688 50.389 68.734 57.179 ;
        RECT 61.926 57.151 68.688 57.225 ;
        RECT 65.238 53.839 72.002 53.911 ;
        RECT 68.642 50.435 68.688 57.225 ;
        RECT 61.88 57.197 68.642 57.271 ;
        RECT 65.284 53.793 72.048 53.865 ;
        RECT 68.596 50.481 68.642 57.271 ;
        RECT 61.834 57.243 68.596 57.317 ;
        RECT 65.33 53.747 72.094 53.819 ;
        RECT 68.55 50.527 68.596 57.317 ;
        RECT 61.788 57.289 68.55 57.363 ;
        RECT 65.376 53.701 72.14 53.773 ;
        RECT 68.504 50.573 68.55 57.363 ;
        RECT 61.742 57.335 68.504 57.409 ;
        RECT 65.422 53.655 72.186 53.727 ;
        RECT 68.458 50.619 68.504 57.409 ;
        RECT 61.696 57.381 68.458 57.455 ;
        RECT 65.468 53.609 72.232 53.681 ;
        RECT 68.412 50.665 68.458 57.455 ;
        RECT 61.65 57.427 68.412 57.501 ;
        RECT 65.514 53.563 72.278 53.635 ;
        RECT 68.366 50.711 68.412 57.501 ;
        RECT 61.604 57.473 68.366 57.547 ;
        RECT 65.56 53.517 80 53.6 ;
        RECT 68.32 50.757 68.366 57.547 ;
        RECT 61.558 57.519 68.32 57.593 ;
        RECT 65.606 53.471 80 53.6 ;
        RECT 68.274 50.803 68.32 57.593 ;
        RECT 61.512 57.565 68.274 57.639 ;
        RECT 65.652 53.425 80 53.6 ;
        RECT 68.228 50.849 68.274 57.639 ;
        RECT 61.466 57.611 68.228 57.685 ;
        RECT 65.698 53.379 80 53.6 ;
        RECT 68.182 50.895 68.228 57.685 ;
        RECT 61.42 57.657 68.182 57.731 ;
        RECT 65.744 53.333 80 53.6 ;
        RECT 68.136 50.941 68.182 57.731 ;
        RECT 61.374 57.703 68.136 57.777 ;
        RECT 65.79 53.287 80 53.6 ;
        RECT 68.09 50.987 68.136 57.777 ;
        RECT 61.328 57.749 68.09 57.823 ;
        RECT 65.836 53.241 80 53.6 ;
        RECT 68.044 51.033 68.09 57.823 ;
        RECT 61.282 57.795 68.044 57.869 ;
        RECT 65.882 53.195 80 53.6 ;
        RECT 67.998 51.079 68.044 57.869 ;
        RECT 61.236 57.841 67.998 57.915 ;
        RECT 65.928 53.149 80 53.6 ;
        RECT 67.952 51.125 67.998 57.915 ;
        RECT 61.19 57.887 67.952 57.961 ;
        RECT 65.974 53.103 80 53.6 ;
        RECT 67.906 51.171 67.952 57.961 ;
        RECT 61.144 57.933 67.906 58.007 ;
        RECT 66.02 53.057 80 53.6 ;
        RECT 67.86 51.217 67.906 58.007 ;
        RECT 61.098 57.979 67.86 58.053 ;
        RECT 66.066 53.011 80 53.6 ;
        RECT 67.814 51.263 67.86 58.053 ;
        RECT 61.052 58.025 67.814 58.099 ;
        RECT 66.112 52.965 80 53.6 ;
        RECT 67.768 51.309 67.814 58.099 ;
        RECT 61.006 58.071 67.768 58.145 ;
        RECT 66.158 52.919 80 53.6 ;
        RECT 67.722 51.355 67.768 58.145 ;
        RECT 60.96 58.117 67.722 58.191 ;
        RECT 66.204 52.873 80 53.6 ;
        RECT 67.676 51.401 67.722 58.191 ;
        RECT 60.914 58.163 67.676 58.237 ;
        RECT 66.25 52.827 80 53.6 ;
        RECT 67.63 51.447 67.676 58.237 ;
        RECT 60.868 58.209 67.63 58.283 ;
        RECT 66.296 52.781 80 53.6 ;
        RECT 67.584 51.493 67.63 58.283 ;
        RECT 60.822 58.255 67.584 58.329 ;
        RECT 66.342 52.735 80 53.6 ;
        RECT 67.538 51.539 67.584 58.329 ;
        RECT 60.776 58.301 67.538 58.375 ;
        RECT 66.388 52.689 80 53.6 ;
        RECT 67.492 51.585 67.538 58.375 ;
        RECT 60.73 58.347 67.492 58.421 ;
        RECT 66.434 52.643 80 53.6 ;
        RECT 67.446 51.631 67.492 58.421 ;
        RECT 60.684 58.393 67.446 58.467 ;
        RECT 66.48 52.597 80 53.6 ;
        RECT 67.4 51.677 67.446 58.467 ;
        RECT 60.638 58.439 67.4 58.513 ;
        RECT 66.526 52.551 80 53.6 ;
        RECT 67.354 51.723 67.4 58.513 ;
        RECT 60.592 58.485 67.354 58.559 ;
        RECT 66.572 52.505 80 53.6 ;
        RECT 67.308 51.769 67.354 58.559 ;
        RECT 60.546 58.531 67.308 58.605 ;
        RECT 66.618 52.459 80 53.6 ;
        RECT 67.262 51.815 67.308 58.605 ;
        RECT 60.5 58.577 67.262 58.651 ;
        RECT 66.664 52.413 80 53.6 ;
        RECT 67.216 51.861 67.262 58.651 ;
        RECT 60.454 58.623 67.216 58.697 ;
        RECT 66.71 52.367 80 53.6 ;
        RECT 67.17 51.907 67.216 58.697 ;
        RECT 60.408 58.669 67.17 58.743 ;
        RECT 66.756 52.321 80 53.6 ;
        RECT 67.124 51.953 67.17 58.743 ;
        RECT 60.362 58.715 67.124 58.789 ;
        RECT 66.802 52.275 80 53.6 ;
        RECT 67.078 51.999 67.124 58.789 ;
        RECT 60.316 58.761 67.078 58.835 ;
        RECT 66.848 52.229 80 53.6 ;
        RECT 67.032 52.045 67.078 58.835 ;
        RECT 60.27 58.807 67.032 58.881 ;
        RECT 66.894 52.183 80 53.6 ;
        RECT 66.986 52.091 67.032 58.881 ;
        RECT 60.224 58.853 66.986 58.927 ;
        RECT 66.94 52.137 80 53.6 ;
        RECT 60.178 58.899 66.94 58.973 ;
        RECT 60.132 58.945 66.894 59.019 ;
        RECT 60.086 58.991 66.848 59.065 ;
        RECT 60.04 59.037 66.802 59.111 ;
        RECT 59.994 59.083 66.756 59.157 ;
        RECT 59.948 59.129 66.71 59.203 ;
        RECT 59.902 59.175 66.664 59.249 ;
        RECT 59.856 59.221 66.618 59.295 ;
        RECT 59.81 59.267 66.572 59.341 ;
        RECT 59.764 59.313 66.526 59.387 ;
        RECT 59.718 59.359 66.48 59.433 ;
        RECT 59.672 59.405 66.434 59.479 ;
        RECT 59.626 59.451 66.388 59.525 ;
        RECT 59.58 59.497 66.342 59.571 ;
        RECT 59.534 59.543 66.296 59.617 ;
        RECT 59.488 59.589 66.25 59.663 ;
        RECT 59.442 59.635 66.204 59.709 ;
        RECT 59.396 59.681 66.158 59.755 ;
        RECT 59.35 59.727 66.112 59.801 ;
        RECT 59.304 59.773 66.066 59.847 ;
        RECT 59.258 59.819 66.02 59.893 ;
        RECT 59.212 59.865 65.974 59.939 ;
        RECT 59.166 59.911 65.928 59.985 ;
        RECT 59.12 59.957 65.882 60.031 ;
        RECT 59.074 60.003 65.836 60.077 ;
        RECT 59.028 60.049 65.79 60.123 ;
        RECT 58.982 60.095 65.744 60.169 ;
        RECT 58.936 60.141 65.698 60.215 ;
        RECT 58.89 60.187 65.652 60.261 ;
        RECT 58.844 60.233 65.606 60.307 ;
        RECT 58.798 60.279 65.56 60.353 ;
        RECT 58.752 60.325 65.514 60.399 ;
        RECT 58.706 60.371 65.468 60.445 ;
        RECT 58.66 60.417 65.422 60.491 ;
        RECT 58.614 60.463 65.376 60.537 ;
        RECT 58.568 60.509 65.33 60.583 ;
        RECT 58.522 60.555 65.284 60.629 ;
        RECT 58.476 60.601 65.238 60.675 ;
        RECT 58.43 60.647 65.192 60.721 ;
        RECT 58.384 60.693 65.146 60.767 ;
        RECT 58.338 60.739 65.1 60.813 ;
        RECT 58.292 60.785 65.054 60.859 ;
        RECT 58.246 60.831 65.008 60.905 ;
        RECT 58.2 60.877 64.962 60.951 ;
        RECT 58.154 60.923 64.916 60.997 ;
        RECT 58.108 60.969 64.87 61.043 ;
        RECT 58.062 61.015 64.824 61.089 ;
        RECT 58.016 61.061 64.778 61.135 ;
        RECT 57.97 61.107 64.732 61.181 ;
        RECT 57.924 61.153 64.686 61.227 ;
        RECT 57.878 61.199 64.64 61.273 ;
        RECT 57.832 61.245 64.594 61.319 ;
        RECT 57.786 61.291 64.548 61.365 ;
        RECT 57.74 61.337 64.502 61.411 ;
        RECT 57.694 61.383 64.456 61.457 ;
        RECT 57.648 61.429 64.41 61.503 ;
        RECT 57.602 61.475 64.364 61.549 ;
        RECT 57.556 61.521 64.318 61.595 ;
        RECT 57.51 61.567 64.272 61.641 ;
        RECT 57.464 61.613 64.226 61.687 ;
        RECT 57.418 61.659 64.18 61.733 ;
        RECT 57.372 61.705 64.134 61.779 ;
        RECT 57.326 61.751 64.088 61.825 ;
        RECT 57.28 61.797 64.042 61.871 ;
        RECT 57.234 61.843 63.996 61.917 ;
        RECT 57.188 61.889 63.95 61.963 ;
        RECT 57.142 61.935 63.904 62.009 ;
        RECT 57.096 61.981 63.858 62.055 ;
        RECT 57.05 62.027 63.812 62.101 ;
        RECT 57.004 62.073 63.766 62.147 ;
        RECT 56.958 62.119 63.72 62.193 ;
        RECT 56.912 62.165 63.674 62.239 ;
        RECT 56.866 62.211 63.628 62.285 ;
        RECT 56.82 62.257 63.582 62.331 ;
        RECT 56.774 62.303 63.536 62.377 ;
        RECT 56.728 62.349 63.49 62.423 ;
        RECT 56.682 62.395 63.444 62.469 ;
        RECT 56.636 62.441 63.398 62.515 ;
        RECT 56.59 62.487 63.352 62.561 ;
        RECT 56.544 62.533 63.306 62.607 ;
        RECT 56.498 62.579 63.26 62.653 ;
        RECT 56.452 62.625 63.214 62.699 ;
        RECT 56.406 62.671 63.168 62.745 ;
        RECT 56.36 62.717 63.122 62.791 ;
        RECT 56.314 62.763 63.076 62.837 ;
        RECT 56.268 62.809 63.03 62.883 ;
        RECT 56.222 62.855 62.984 62.929 ;
        RECT 56.176 62.901 62.938 62.975 ;
        RECT 56.13 62.947 62.892 63.021 ;
        RECT 56.084 62.993 62.846 63.067 ;
        RECT 56.038 63.039 62.8 63.113 ;
        RECT 55.992 63.085 62.754 63.159 ;
        RECT 55.946 63.131 62.708 63.205 ;
        RECT 55.9 63.177 62.662 63.251 ;
        RECT 55.854 63.223 62.616 63.297 ;
        RECT 55.808 63.269 62.57 63.343 ;
        RECT 55.762 63.315 62.524 63.389 ;
        RECT 55.716 63.361 62.478 63.435 ;
        RECT 55.67 63.407 62.432 63.481 ;
        RECT 55.624 63.453 62.386 63.527 ;
        RECT 55.578 63.499 62.34 63.573 ;
        RECT 55.532 63.545 62.294 63.619 ;
        RECT 55.486 63.591 62.248 63.665 ;
        RECT 55.44 63.637 62.202 63.711 ;
        RECT 55.394 63.683 62.156 63.757 ;
        RECT 55.348 63.729 62.11 63.803 ;
        RECT 55.302 63.775 62.064 63.849 ;
        RECT 55.256 63.821 62.018 63.895 ;
        RECT 55.21 63.867 61.972 63.941 ;
        RECT 55.164 63.913 61.926 63.987 ;
        RECT 55.118 63.959 61.88 64.033 ;
        RECT 55.072 64.005 61.834 64.079 ;
        RECT 55.026 64.051 61.788 64.125 ;
        RECT 54.98 64.097 61.742 64.171 ;
        RECT 54.934 64.143 61.696 64.217 ;
        RECT 54.888 64.189 61.65 64.263 ;
        RECT 54.842 64.235 61.604 64.309 ;
        RECT 54.796 64.281 61.558 64.355 ;
        RECT 54.75 64.327 61.512 64.401 ;
        RECT 54.704 64.373 61.466 64.447 ;
        RECT 54.658 64.419 61.42 64.493 ;
        RECT 54.612 64.465 61.374 64.539 ;
        RECT 54.566 64.511 61.328 64.585 ;
        RECT 54.52 64.557 61.282 64.631 ;
        RECT 54.474 64.603 61.236 64.677 ;
        RECT 54.428 64.649 61.19 64.723 ;
        RECT 54.382 64.695 61.144 64.769 ;
        RECT 54.336 64.741 61.098 64.815 ;
        RECT 54.29 64.787 61.052 64.861 ;
        RECT 54.244 64.833 61.006 64.907 ;
        RECT 54.198 64.879 60.96 64.953 ;
        RECT 54.152 64.925 60.914 64.999 ;
        RECT 54.106 64.971 60.868 65.045 ;
        RECT 54.06 65.017 60.822 65.091 ;
        RECT 54.014 65.063 60.776 65.137 ;
        RECT 53.968 65.109 60.73 65.183 ;
        RECT 53.922 65.155 60.684 65.229 ;
        RECT 53.876 65.201 60.638 65.275 ;
        RECT 53.83 65.247 60.592 65.321 ;
        RECT 53.784 65.293 60.546 65.367 ;
        RECT 53.738 65.339 60.5 65.413 ;
        RECT 53.692 65.385 60.454 65.459 ;
        RECT 53.646 65.431 60.408 65.505 ;
        RECT 53.584 65.508 60.362 65.551 ;
        RECT 53.6 65.477 60.362 65.551 ;
        RECT 53.538 65.539 60.316 65.597 ;
        RECT 53.492 65.585 60.27 65.643 ;
        RECT 53.446 65.631 60.224 65.689 ;
        RECT 53.4 65.677 60.178 65.735 ;
        RECT 53.354 65.723 60.132 65.781 ;
        RECT 53.308 65.769 60.086 65.827 ;
        RECT 53.262 65.815 60.04 65.873 ;
        RECT 53.216 65.861 59.994 65.919 ;
        RECT 53.17 65.907 59.948 65.965 ;
        RECT 53.124 65.953 59.902 66.011 ;
        RECT 53.078 65.999 59.856 66.057 ;
        RECT 53.032 66.045 59.81 66.103 ;
        RECT 52.986 66.091 59.764 66.149 ;
        RECT 52.94 66.137 59.718 66.195 ;
        RECT 52.894 66.183 59.672 66.241 ;
        RECT 52.848 66.229 59.626 66.287 ;
        RECT 52.802 66.275 59.58 66.333 ;
        RECT 52.756 66.321 59.534 66.379 ;
        RECT 52.71 66.367 59.488 66.425 ;
        RECT 52.664 66.413 59.442 66.471 ;
        RECT 52.618 66.459 59.396 66.517 ;
        RECT 52.572 66.505 59.35 66.563 ;
        RECT 52.526 66.551 59.304 66.609 ;
        RECT 52.48 66.597 59.258 66.655 ;
        RECT 52.434 66.643 59.212 66.701 ;
        RECT 52.388 66.689 59.166 66.747 ;
        RECT 52.342 66.735 59.12 66.793 ;
        RECT 52.296 66.781 59.074 66.839 ;
        RECT 52.25 66.827 59.028 66.885 ;
        RECT 52.204 66.873 58.982 66.931 ;
        RECT 52.158 66.919 58.936 66.977 ;
        RECT 52.112 66.965 58.89 67.023 ;
        RECT 52.066 67.011 58.844 67.069 ;
        RECT 52.02 67.057 58.798 67.115 ;
        RECT 51.974 67.103 58.752 67.161 ;
        RECT 51.928 67.149 58.706 67.207 ;
        RECT 51.882 67.195 58.66 67.253 ;
        RECT 51.836 67.241 58.614 67.299 ;
        RECT 51.79 67.287 58.568 67.345 ;
        RECT 51.744 67.333 58.522 67.391 ;
        RECT 51.698 67.379 58.476 67.437 ;
        RECT 51.652 67.425 58.43 67.483 ;
        RECT 51.606 67.471 58.384 67.529 ;
        RECT 51.56 67.517 58.338 67.575 ;
        RECT 51.514 67.563 58.292 67.621 ;
        RECT 51.468 67.609 58.246 67.667 ;
        RECT 51.422 67.655 58.2 67.713 ;
        RECT 51.376 67.701 58.154 67.759 ;
        RECT 51.33 67.747 58.108 67.805 ;
        RECT 51.284 67.793 58.062 67.851 ;
        RECT 51.238 67.839 58.016 67.897 ;
        RECT 51.192 67.885 57.97 67.943 ;
        RECT 51.146 67.931 57.924 67.989 ;
        RECT 51.1 67.977 57.878 68.035 ;
        RECT 51.054 68.023 57.832 68.081 ;
        RECT 51.008 68.069 57.786 68.127 ;
        RECT 50.962 68.115 57.74 68.173 ;
        RECT 50.916 68.161 57.694 68.219 ;
        RECT 50.87 68.207 57.648 68.265 ;
        RECT 50.824 68.253 57.602 68.311 ;
        RECT 50.778 68.299 57.556 68.357 ;
        RECT 50.732 68.345 57.51 68.403 ;
        RECT 50.686 68.391 57.464 68.449 ;
        RECT 50.64 68.437 57.418 68.495 ;
        RECT 50.594 68.483 57.372 68.541 ;
        RECT 50.548 68.529 57.326 68.587 ;
        RECT 50.502 68.575 57.28 68.633 ;
        RECT 50.456 68.621 57.234 68.679 ;
        RECT 50.41 68.667 57.188 68.725 ;
        RECT 50.364 68.713 57.142 68.771 ;
        RECT 50.318 68.759 57.096 68.817 ;
        RECT 50.272 68.805 57.05 68.863 ;
        RECT 50.226 68.851 57.004 68.909 ;
        RECT 50.18 68.897 56.958 68.955 ;
        RECT 50.134 68.943 56.912 69.001 ;
        RECT 50.088 68.989 56.866 69.047 ;
        RECT 50.042 69.035 56.82 69.093 ;
        RECT 49.996 69.081 56.774 69.139 ;
        RECT 49.95 69.127 56.728 69.185 ;
        RECT 49.904 69.173 56.682 69.231 ;
        RECT 49.858 69.219 56.636 69.277 ;
        RECT 49.812 69.265 56.59 69.323 ;
        RECT 49.766 69.311 56.544 69.369 ;
        RECT 49.72 69.357 56.498 69.415 ;
        RECT 49.674 69.403 56.452 69.461 ;
        RECT 49.628 69.449 56.406 69.507 ;
        RECT 49.582 69.495 56.36 69.553 ;
        RECT 49.536 69.541 56.314 69.599 ;
        RECT 49.49 69.587 56.268 69.645 ;
        RECT 49.444 69.633 56.222 69.691 ;
        RECT 49.398 69.679 56.176 69.737 ;
        RECT 49.352 69.725 56.13 69.783 ;
        RECT 49.306 69.771 56.084 69.829 ;
        RECT 49.26 69.817 56.038 69.875 ;
        RECT 49.214 69.863 55.992 69.921 ;
        RECT 49.168 69.909 55.946 69.967 ;
        RECT 49.122 69.955 55.9 70.013 ;
        RECT 49.076 70.001 55.854 70.059 ;
        RECT 49.03 70.047 55.808 70.105 ;
        RECT 48.984 70.093 55.762 70.151 ;
        RECT 48.938 70.139 55.716 70.197 ;
        RECT 48.892 70.185 55.67 70.243 ;
        RECT 48.846 70.231 55.624 70.289 ;
        RECT 48.8 70.277 55.578 70.335 ;
        RECT 48.8 70.277 55.532 70.381 ;
        RECT 48.8 70.277 55.486 70.427 ;
        RECT 48.8 70.277 55.44 70.473 ;
        RECT 48.8 70.277 55.394 70.519 ;
        RECT 48.8 70.277 55.348 70.565 ;
        RECT 48.8 70.277 55.302 70.611 ;
        RECT 48.8 70.277 55.256 70.657 ;
        RECT 48.8 70.277 55.21 70.703 ;
        RECT 48.8 70.277 55.164 70.749 ;
        RECT 48.8 70.277 55.118 70.795 ;
        RECT 48.8 70.277 55.072 70.841 ;
        RECT 48.8 70.277 55.026 70.887 ;
        RECT 48.8 70.277 54.98 70.933 ;
        RECT 48.8 70.277 54.934 70.979 ;
        RECT 48.8 70.277 54.888 71.025 ;
        RECT 48.8 70.277 54.842 71.071 ;
        RECT 48.8 70.277 54.796 71.117 ;
        RECT 48.8 70.277 54.75 71.163 ;
        RECT 48.8 70.277 54.704 71.209 ;
        RECT 48.8 70.277 54.658 71.255 ;
        RECT 48.8 70.277 54.612 71.301 ;
        RECT 48.8 70.277 54.566 71.347 ;
        RECT 48.8 70.277 54.52 71.393 ;
        RECT 48.8 70.277 54.474 71.439 ;
        RECT 48.8 70.277 54.428 71.485 ;
        RECT 48.8 70.277 54.382 71.531 ;
        RECT 48.8 70.277 54.336 71.577 ;
        RECT 48.8 70.277 54.29 71.623 ;
        RECT 48.8 70.277 54.244 71.669 ;
        RECT 48.8 70.277 54.198 71.715 ;
        RECT 48.8 70.277 54.152 71.761 ;
        RECT 48.8 70.277 54.106 71.807 ;
        RECT 48.8 70.277 54.06 71.853 ;
        RECT 48.8 70.277 54.014 71.899 ;
        RECT 48.8 70.277 53.968 71.945 ;
        RECT 48.8 70.277 53.922 71.991 ;
        RECT 48.8 70.277 53.876 72.037 ;
        RECT 48.8 70.277 53.83 72.083 ;
        RECT 48.8 70.277 53.784 72.129 ;
        RECT 48.8 70.277 53.738 72.175 ;
        RECT 48.8 70.277 53.692 72.221 ;
        RECT 48.8 70.277 53.646 72.267 ;
        RECT 48.8 70.277 53.6 80 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 80 ;
    LAYER M1 ;
      RECT 0 0 80 80 ;
    LAYER V1 ;
      RECT 0 0 80 80 ;
    LAYER M2 ;
      RECT 0 0 80 80 ;
    LAYER A1 ;
      RECT 0 0 80 80 ;
    LAYER C2 ;
      RECT 0 0 80 80 ;
    LAYER CB ;
      RECT 0 0 80 80 ;
    LAYER JV ;
      RECT 0 0 80 80 ;
    LAYER YS ;
      RECT 0 0 80 80 ;
    LAYER JW ;
      RECT 0 0 80 80 ;
    LAYER QB ;
      RECT 0 0 80 80 ;
    LAYER QA ;
      RECT 0 0 80 80 ;
    LAYER JA ;
      RECT 0 0 80 80 ;
    LAYER AY ;
      RECT 0 0 80 80 ;
    LAYER C1 ;
      RECT 0 0 80 80 ;
    LAYER C5 ;
      RECT 0 0 80 80 ;
    LAYER C4 ;
      RECT 0 0 80 80 ;
    LAYER C3 ;
      RECT 0 0 80 80 ;
    LAYER A4 ;
      RECT 0 0 80 80 ;
    LAYER A3 ;
      RECT 0 0 80 80 ;
    LAYER A2 ;
      RECT 0 0 80 80 ;
  END
END RIIO_EG1D80V_CORNER_45

MACRO RIIO_EG1D80V_CORNER_EG
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CORNER_EG 0 0 ;
  SIZE 80 BY 80 ;
  SYMMETRY X Y ;
  SITE corner_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 24 24 78.4 28.8 ;
        RECT 24 24 28.8 78.4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 42.6 80 47.4 ;
        RECT 42.6 42.6 47.4 80 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 17.8 80 22.6 ;
        RECT 17.8 17.8 22.6 80 ;
    END
    PORT
      LAYER QB ;
        RECT 5.4 5.4 80 10.2 ;
        RECT 5.4 5.4 10.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 0 73.6 2.4 78.4 ;
      LAYER JA ;
        RECT 0 73.6 2.4 78.4 ;
      LAYER QB ;
        RECT 0 73.6 2.4 78.4 ;
    END
    PORT
      LAYER QA ;
        RECT 0 67.4 2.4 72.2 ;
      LAYER JA ;
        RECT 0 67.4 2.4 72.2 ;
      LAYER QB ;
        RECT 0 67.4 2.4 72.2 ;
    END
    PORT
      LAYER QA ;
        RECT 0 61.2 2.4 66 ;
      LAYER JA ;
        RECT 0 61.2 2.4 66 ;
      LAYER QB ;
        RECT 0 61.2 2.4 66 ;
    END
    PORT
      LAYER QA ;
        RECT 0 55 2.4 59.8 ;
      LAYER JA ;
        RECT 0 55 2.4 59.8 ;
      LAYER QB ;
        RECT 0 55 2.4 59.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 48.8 2.4 53.6 ;
      LAYER JA ;
        RECT 0 48.8 2.4 53.6 ;
      LAYER QB ;
        RECT 0 48.8 2.4 53.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 42.6 2.4 47.4 ;
      LAYER JA ;
        RECT 0 42.6 2.4 47.4 ;
      LAYER QB ;
        RECT 0 42.6 2.4 47.4 ;
    END
    PORT
      LAYER QA ;
        RECT 0 36.4 2.4 41.2 ;
      LAYER JA ;
        RECT 0 36.4 2.4 41.2 ;
      LAYER QB ;
        RECT 0 36.4 2.4 41.2 ;
    END
    PORT
      LAYER QA ;
        RECT 0 30.2 2.4 35 ;
      LAYER JA ;
        RECT 0 30.2 2.4 35 ;
      LAYER QB ;
        RECT 0 30.2 2.4 35 ;
    END
    PORT
      LAYER QA ;
        RECT 0 24 2.4 28.8 ;
      LAYER JA ;
        RECT 0 24 2.4 28.8 ;
      LAYER QB ;
        RECT 0 24 2.4 28.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 17.8 2.4 22.6 ;
      LAYER JA ;
        RECT 0 17.8 2.4 22.6 ;
      LAYER QB ;
        RECT 0 17.8 2.4 22.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 11.6 2.4 16.4 ;
      LAYER JA ;
        RECT 0 11.6 2.4 16.4 ;
      LAYER QB ;
        RECT 0 11.6 2.4 16.4 ;
    END
    PORT
      LAYER QA ;
        RECT 0 5.4 2.4 10.2 ;
      LAYER JA ;
        RECT 0 5.4 2.4 10.2 ;
      LAYER QB ;
        RECT 0 5.4 2.4 10.2 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 36.4 36.4 80 41.2 ;
        RECT 36.4 36.4 41.2 80 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 30.2 80 35 ;
        RECT 30.2 30.2 35 80 ;
    END
    PORT
      LAYER QB ;
        RECT 11.6 11.6 80 16.4 ;
        RECT 11.6 11.6 16.4 80 ;
    END
    PORT
      LAYER QA ;
        RECT 5.4 0 10.2 2.4 ;
      LAYER JA ;
        RECT 5.4 0 10.2 2.4 ;
      LAYER QB ;
        RECT 5.4 0 10.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 11.6 0 16.4 2.4 ;
      LAYER JA ;
        RECT 11.6 0 16.4 2.4 ;
      LAYER QB ;
        RECT 11.6 0 16.4 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 17.8 0 22.6 2.4 ;
      LAYER JA ;
        RECT 17.8 0 22.6 2.4 ;
      LAYER QB ;
        RECT 17.8 0 22.6 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 24 0 28.8 2.4 ;
      LAYER JA ;
        RECT 24 0 28.8 2.4 ;
      LAYER QB ;
        RECT 24 0 28.8 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 30.2 0 35 2.4 ;
      LAYER JA ;
        RECT 30.2 0 35 2.4 ;
      LAYER QB ;
        RECT 30.2 0 35 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 36.4 0 41.2 2.4 ;
      LAYER JA ;
        RECT 36.4 0 41.2 2.4 ;
      LAYER QB ;
        RECT 36.4 0 41.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 42.6 0 47.4 2.4 ;
      LAYER JA ;
        RECT 42.6 0 47.4 2.4 ;
      LAYER QB ;
        RECT 42.6 0 47.4 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 48.8 0 53.6 2.4 ;
      LAYER JA ;
        RECT 48.8 0 53.6 2.4 ;
      LAYER QB ;
        RECT 48.8 0 53.6 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 55 0 59.8 2.4 ;
      LAYER JA ;
        RECT 55 0 59.8 2.4 ;
      LAYER QB ;
        RECT 55 0 59.8 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 61.2 0 66 2.4 ;
      LAYER JA ;
        RECT 61.2 0 66 2.4 ;
      LAYER QB ;
        RECT 61.2 0 66 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 67.4 0 72.2 2.4 ;
      LAYER JA ;
        RECT 67.4 0 72.2 2.4 ;
      LAYER QB ;
        RECT 67.4 0 72.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 73.6 0 78.4 2.4 ;
      LAYER JA ;
        RECT 73.6 0 78.4 2.4 ;
      LAYER QB ;
        RECT 73.6 0 78.4 2.4 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 61.2 61.2 80 66 ;
        RECT 61.2 61.2 66 80 ;
    END
    PORT
      LAYER QB ;
        RECT 55 55 80 59.8 ;
        RECT 55 55 59.8 80 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 67.4 67.4 80 72.2 ;
        RECT 67.4 67.4 72.2 80 ;
    END
    PORT
      LAYER QB ;
        RECT 48.8 48.8 80 53.6 ;
        RECT 48.8 48.8 53.6 80 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 80 ;
    LAYER M1 ;
      RECT 0 0 80 80 ;
    LAYER V1 ;
      RECT 0 0 80 80 ;
    LAYER M2 ;
      RECT 0 0 80 80 ;
    LAYER A1 ;
      RECT 0 0 80 80 ;
    LAYER C2 ;
      RECT 0 0 80 80 ;
    LAYER CB ;
      RECT 0 0 80 80 ;
    LAYER JV ;
      RECT 0 0 80 80 ;
    LAYER YS ;
      RECT 0 0 80 80 ;
    LAYER JW ;
      RECT 0 0 80 80 ;
    LAYER QB ;
      RECT 0 0 80 80 ;
    LAYER QA ;
      RECT 0 0 80 80 ;
    LAYER JA ;
      RECT 0 0 80 80 ;
    LAYER AY ;
      RECT 0 0 80 80 ;
    LAYER C1 ;
      RECT 0 0 80 80 ;
    LAYER C5 ;
      RECT 0 0 80 80 ;
    LAYER C4 ;
      RECT 0 0 80 80 ;
    LAYER C3 ;
      RECT 0 0 80 80 ;
    LAYER A4 ;
      RECT 0 0 80 80 ;
    LAYER A3 ;
      RECT 0 0 80 80 ;
    LAYER A2 ;
      RECT 0 0 80 80 ;
  END
END RIIO_EG1D80V_CORNER_EG

MACRO RIIO_EG1D80V_CORNER_HVT
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CORNER_HVT 0 0 ;
  SIZE 80 BY 80 ;
  SYMMETRY X Y ;
  SITE corner_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 67.4 67.4 80 72.2 ;
        RECT 67.4 67.4 72.2 80 ;
    END
    PORT
      LAYER QB ;
        RECT 48.8 48.8 80 53.6 ;
        RECT 48.8 48.8 53.6 80 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 24 24 78.4 28.8 ;
        RECT 24 24 28.8 78.4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 42.6 80 47.4 ;
        RECT 42.6 42.6 47.4 80 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 17.8 80 22.6 ;
        RECT 17.8 17.8 22.6 80 ;
    END
    PORT
      LAYER QB ;
        RECT 5.4 5.4 80 10.2 ;
        RECT 5.4 5.4 10.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 0 73.6 2.4 78.4 ;
      LAYER JA ;
        RECT 0 73.6 2.4 78.4 ;
      LAYER QB ;
        RECT 0 73.6 2.4 78.4 ;
    END
    PORT
      LAYER QA ;
        RECT 0 67.4 2.4 72.2 ;
      LAYER JA ;
        RECT 0 67.4 2.4 72.2 ;
      LAYER QB ;
        RECT 0 67.4 2.4 72.2 ;
    END
    PORT
      LAYER QA ;
        RECT 0 61.2 2.4 66 ;
      LAYER JA ;
        RECT 0 61.2 2.4 66 ;
      LAYER QB ;
        RECT 0 61.2 2.4 66 ;
    END
    PORT
      LAYER QA ;
        RECT 0 55 2.4 59.8 ;
      LAYER JA ;
        RECT 0 55 2.4 59.8 ;
      LAYER QB ;
        RECT 0 55 2.4 59.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 48.8 2.4 53.6 ;
      LAYER JA ;
        RECT 0 48.8 2.4 53.6 ;
      LAYER QB ;
        RECT 0 48.8 2.4 53.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 42.6 2.4 47.4 ;
      LAYER JA ;
        RECT 0 42.6 2.4 47.4 ;
      LAYER QB ;
        RECT 0 42.6 2.4 47.4 ;
    END
    PORT
      LAYER QA ;
        RECT 0 36.4 2.4 41.2 ;
      LAYER JA ;
        RECT 0 36.4 2.4 41.2 ;
      LAYER QB ;
        RECT 0 36.4 2.4 41.2 ;
    END
    PORT
      LAYER QA ;
        RECT 0 30.2 2.4 35 ;
      LAYER JA ;
        RECT 0 30.2 2.4 35 ;
      LAYER QB ;
        RECT 0 30.2 2.4 35 ;
    END
    PORT
      LAYER QA ;
        RECT 0 24 2.4 28.8 ;
      LAYER JA ;
        RECT 0 24 2.4 28.8 ;
      LAYER QB ;
        RECT 0 24 2.4 28.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 17.8 2.4 22.6 ;
      LAYER JA ;
        RECT 0 17.8 2.4 22.6 ;
      LAYER QB ;
        RECT 0 17.8 2.4 22.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 11.6 2.4 16.4 ;
      LAYER JA ;
        RECT 0 11.6 2.4 16.4 ;
      LAYER QB ;
        RECT 0 11.6 2.4 16.4 ;
    END
    PORT
      LAYER QA ;
        RECT 0 5.4 2.4 10.2 ;
      LAYER JA ;
        RECT 0 5.4 2.4 10.2 ;
      LAYER QB ;
        RECT 0 5.4 2.4 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 61.2 61.2 80 66 ;
        RECT 61.2 61.2 66 80 ;
    END
    PORT
      LAYER QB ;
        RECT 55 55 80 59.8 ;
        RECT 55 55 59.8 80 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 36.4 36.4 80 41.2 ;
        RECT 36.4 36.4 41.2 80 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 30.2 80 35 ;
        RECT 30.2 30.2 35 80 ;
    END
    PORT
      LAYER QB ;
        RECT 11.6 11.6 80 16.4 ;
        RECT 11.6 11.6 16.4 80 ;
    END
    PORT
      LAYER QA ;
        RECT 5.4 0 10.2 2.4 ;
      LAYER JA ;
        RECT 5.4 0 10.2 2.4 ;
      LAYER QB ;
        RECT 5.4 0 10.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 11.6 0 16.4 2.4 ;
      LAYER JA ;
        RECT 11.6 0 16.4 2.4 ;
      LAYER QB ;
        RECT 11.6 0 16.4 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 17.8 0 22.6 2.4 ;
      LAYER JA ;
        RECT 17.8 0 22.6 2.4 ;
      LAYER QB ;
        RECT 17.8 0 22.6 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 24 0 28.8 2.4 ;
      LAYER JA ;
        RECT 24 0 28.8 2.4 ;
      LAYER QB ;
        RECT 24 0 28.8 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 30.2 0 35 2.4 ;
      LAYER JA ;
        RECT 30.2 0 35 2.4 ;
      LAYER QB ;
        RECT 30.2 0 35 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 36.4 0 41.2 2.4 ;
      LAYER JA ;
        RECT 36.4 0 41.2 2.4 ;
      LAYER QB ;
        RECT 36.4 0 41.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 42.6 0 47.4 2.4 ;
      LAYER JA ;
        RECT 42.6 0 47.4 2.4 ;
      LAYER QB ;
        RECT 42.6 0 47.4 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 48.8 0 53.6 2.4 ;
      LAYER JA ;
        RECT 48.8 0 53.6 2.4 ;
      LAYER QB ;
        RECT 48.8 0 53.6 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 55 0 59.8 2.4 ;
      LAYER JA ;
        RECT 55 0 59.8 2.4 ;
      LAYER QB ;
        RECT 55 0 59.8 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 61.2 0 66 2.4 ;
      LAYER JA ;
        RECT 61.2 0 66 2.4 ;
      LAYER QB ;
        RECT 61.2 0 66 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 67.4 0 72.2 2.4 ;
      LAYER JA ;
        RECT 67.4 0 72.2 2.4 ;
      LAYER QB ;
        RECT 67.4 0 72.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 73.6 0 78.4 2.4 ;
      LAYER JA ;
        RECT 73.6 0 78.4 2.4 ;
      LAYER QB ;
        RECT 73.6 0 78.4 2.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 80 ;
    LAYER M1 ;
      RECT 0 0 80 80 ;
    LAYER V1 ;
      RECT 0 0 80 80 ;
    LAYER M2 ;
      RECT 0 0 80 80 ;
    LAYER A1 ;
      RECT 0 0 80 80 ;
    LAYER C2 ;
      RECT 0 0 80 80 ;
    LAYER CB ;
      RECT 0 0 80 80 ;
    LAYER JV ;
      RECT 0 0 80 80 ;
    LAYER YS ;
      RECT 0 0 80 80 ;
    LAYER JW ;
      RECT 0 0 80 80 ;
    LAYER QB ;
      RECT 0 0 80 80 ;
    LAYER QA ;
      RECT 0 0 80 80 ;
    LAYER JA ;
      RECT 0 0 80 80 ;
    LAYER AY ;
      RECT 0 0 80 80 ;
    LAYER C1 ;
      RECT 0 0 80 80 ;
    LAYER C5 ;
      RECT 0 0 80 80 ;
    LAYER C4 ;
      RECT 0 0 80 80 ;
    LAYER C3 ;
      RECT 0 0 80 80 ;
    LAYER A4 ;
      RECT 0 0 80 80 ;
    LAYER A3 ;
      RECT 0 0 80 80 ;
    LAYER A2 ;
      RECT 0 0 80 80 ;
  END
END RIIO_EG1D80V_CORNER_HVT

MACRO RIIO_EG1D80V_CORNER_RVT
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CORNER_RVT 0 0 ;
  SIZE 80 BY 80 ;
  SYMMETRY X Y ;
  SITE corner_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 67.4 67.4 80 72.2 ;
        RECT 67.4 67.4 72.2 80 ;
    END
    PORT
      LAYER QB ;
        RECT 48.8 48.8 80 53.6 ;
        RECT 48.8 48.8 53.6 80 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 61.2 61.2 80 66 ;
        RECT 61.2 61.2 66 80 ;
    END
    PORT
      LAYER QB ;
        RECT 55 55 80 59.8 ;
        RECT 55 55 59.8 80 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 36.4 36.4 80 41.2 ;
        RECT 36.4 36.4 41.2 80 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 30.2 80 35 ;
        RECT 30.2 30.2 35 80 ;
    END
    PORT
      LAYER QB ;
        RECT 11.6 11.6 80 16.4 ;
        RECT 11.6 11.6 16.4 80 ;
    END
    PORT
      LAYER QA ;
        RECT 5.4 0 10.2 2.4 ;
      LAYER JA ;
        RECT 5.4 0 10.2 2.4 ;
      LAYER QB ;
        RECT 5.4 0 10.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 11.6 0 16.4 2.4 ;
      LAYER JA ;
        RECT 11.6 0 16.4 2.4 ;
      LAYER QB ;
        RECT 11.6 0 16.4 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 17.8 0 22.6 2.4 ;
      LAYER JA ;
        RECT 17.8 0 22.6 2.4 ;
      LAYER QB ;
        RECT 17.8 0 22.6 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 24 0 28.8 2.4 ;
      LAYER JA ;
        RECT 24 0 28.8 2.4 ;
      LAYER QB ;
        RECT 24 0 28.8 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 30.2 0 35 2.4 ;
      LAYER JA ;
        RECT 30.2 0 35 2.4 ;
      LAYER QB ;
        RECT 30.2 0 35 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 36.4 0 41.2 2.4 ;
      LAYER JA ;
        RECT 36.4 0 41.2 2.4 ;
      LAYER QB ;
        RECT 36.4 0 41.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 42.6 0 47.4 2.4 ;
      LAYER JA ;
        RECT 42.6 0 47.4 2.4 ;
      LAYER QB ;
        RECT 42.6 0 47.4 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 48.8 0 53.6 2.4 ;
      LAYER JA ;
        RECT 48.8 0 53.6 2.4 ;
      LAYER QB ;
        RECT 48.8 0 53.6 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 55 0 59.8 2.4 ;
      LAYER JA ;
        RECT 55 0 59.8 2.4 ;
      LAYER QB ;
        RECT 55 0 59.8 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 61.2 0 66 2.4 ;
      LAYER JA ;
        RECT 61.2 0 66 2.4 ;
      LAYER QB ;
        RECT 61.2 0 66 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 67.4 0 72.2 2.4 ;
      LAYER JA ;
        RECT 67.4 0 72.2 2.4 ;
      LAYER QB ;
        RECT 67.4 0 72.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 73.6 0 78.4 2.4 ;
      LAYER JA ;
        RECT 73.6 0 78.4 2.4 ;
      LAYER QB ;
        RECT 73.6 0 78.4 2.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 24 24 78.4 28.8 ;
        RECT 24 24 28.8 78.4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 42.6 80 47.4 ;
        RECT 42.6 42.6 47.4 80 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 17.8 80 22.6 ;
        RECT 17.8 17.8 22.6 80 ;
    END
    PORT
      LAYER QB ;
        RECT 5.4 5.4 80 10.2 ;
        RECT 5.4 5.4 10.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 0 73.6 2.4 78.4 ;
      LAYER JA ;
        RECT 0 73.6 2.4 78.4 ;
      LAYER QB ;
        RECT 0 73.6 2.4 78.4 ;
    END
    PORT
      LAYER QA ;
        RECT 0 67.4 2.4 72.2 ;
      LAYER JA ;
        RECT 0 67.4 2.4 72.2 ;
      LAYER QB ;
        RECT 0 67.4 2.4 72.2 ;
    END
    PORT
      LAYER QA ;
        RECT 0 61.2 2.4 66 ;
      LAYER JA ;
        RECT 0 61.2 2.4 66 ;
      LAYER QB ;
        RECT 0 61.2 2.4 66 ;
    END
    PORT
      LAYER QA ;
        RECT 0 55 2.4 59.8 ;
      LAYER JA ;
        RECT 0 55 2.4 59.8 ;
      LAYER QB ;
        RECT 0 55 2.4 59.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 48.8 2.4 53.6 ;
      LAYER JA ;
        RECT 0 48.8 2.4 53.6 ;
      LAYER QB ;
        RECT 0 48.8 2.4 53.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 42.6 2.4 47.4 ;
      LAYER JA ;
        RECT 0 42.6 2.4 47.4 ;
      LAYER QB ;
        RECT 0 42.6 2.4 47.4 ;
    END
    PORT
      LAYER QA ;
        RECT 0 36.4 2.4 41.2 ;
      LAYER JA ;
        RECT 0 36.4 2.4 41.2 ;
      LAYER QB ;
        RECT 0 36.4 2.4 41.2 ;
    END
    PORT
      LAYER QA ;
        RECT 0 30.2 2.4 35 ;
      LAYER JA ;
        RECT 0 30.2 2.4 35 ;
      LAYER QB ;
        RECT 0 30.2 2.4 35 ;
    END
    PORT
      LAYER QA ;
        RECT 0 24 2.4 28.8 ;
      LAYER JA ;
        RECT 0 24 2.4 28.8 ;
      LAYER QB ;
        RECT 0 24 2.4 28.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 17.8 2.4 22.6 ;
      LAYER JA ;
        RECT 0 17.8 2.4 22.6 ;
      LAYER QB ;
        RECT 0 17.8 2.4 22.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 11.6 2.4 16.4 ;
      LAYER JA ;
        RECT 0 11.6 2.4 16.4 ;
      LAYER QB ;
        RECT 0 11.6 2.4 16.4 ;
    END
    PORT
      LAYER QA ;
        RECT 0 5.4 2.4 10.2 ;
      LAYER JA ;
        RECT 0 5.4 2.4 10.2 ;
      LAYER QB ;
        RECT 0 5.4 2.4 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 80 80 ;
    LAYER M1 ;
      RECT 0 0 80 80 ;
    LAYER V1 ;
      RECT 0 0 80 80 ;
    LAYER M2 ;
      RECT 0 0 80 80 ;
    LAYER A1 ;
      RECT 0 0 80 80 ;
    LAYER C2 ;
      RECT 0 0 80 80 ;
    LAYER CB ;
      RECT 0 0 80 80 ;
    LAYER JV ;
      RECT 0 0 80 80 ;
    LAYER YS ;
      RECT 0 0 80 80 ;
    LAYER JW ;
      RECT 0 0 80 80 ;
    LAYER QB ;
      RECT 0 0 80 80 ;
    LAYER QA ;
      RECT 0 0 80 80 ;
    LAYER JA ;
      RECT 0 0 80 80 ;
    LAYER AY ;
      RECT 0 0 80 80 ;
    LAYER C1 ;
      RECT 0 0 80 80 ;
    LAYER C5 ;
      RECT 0 0 80 80 ;
    LAYER C4 ;
      RECT 0 0 80 80 ;
    LAYER C3 ;
      RECT 0 0 80 80 ;
    LAYER A4 ;
      RECT 0 0 80 80 ;
    LAYER A3 ;
      RECT 0 0 80 80 ;
    LAYER A2 ;
      RECT 0 0 80 80 ;
  END
END RIIO_EG1D80V_CORNER_RVT

MACRO RIIO_EG1D80V_ANACORE_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ANACORE_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VESD3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 63.22955 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 62.855 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 52.45 78.15 52.95 80 ;
        RECT 51.675 78.15 52.175 80 ;
        RECT 50.9 78.15 51.4 80 ;
        RECT 50.125 78.15 50.625 80 ;
        RECT 49.35 78.15 49.85 80 ;
      LAYER M2 ;
        RECT 52.45 78.15 52.95 80 ;
        RECT 51.675 78.15 52.175 80 ;
        RECT 50.9 78.15 51.4 80 ;
        RECT 50.125 78.15 50.625 80 ;
        RECT 49.35 78.15 49.85 80 ;
      LAYER C1 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER JA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER QB ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER QA ;
        RECT 49.65 77.975 52.65 80 ;
    END
  END VESD3_B
  PIN VRES1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 75.6725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 19.55 78.15 20.05 80 ;
        RECT 18.775 78.15 19.275 80 ;
        RECT 18 78.15 18.5 80 ;
        RECT 17.225 78.15 17.725 80 ;
        RECT 16.45 78.15 16.95 80 ;
      LAYER M2 ;
        RECT 19.55 78.15 20.05 80 ;
        RECT 18.775 78.15 19.275 80 ;
        RECT 18 78.15 18.5 80 ;
        RECT 17.225 78.15 17.725 80 ;
        RECT 16.45 78.15 16.95 80 ;
      LAYER C1 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER JA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER QB ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER QA ;
        RECT 16.75 77.975 19.75 80 ;
    END
  END VRES1_B
  PIN VRES0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 72.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 16.735 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.105 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 14.85 78.15 15.35 80 ;
        RECT 14.075 78.15 14.575 80 ;
        RECT 13.3 78.15 13.8 80 ;
        RECT 12.525 78.15 13.025 80 ;
        RECT 11.75 78.15 12.25 80 ;
      LAYER M2 ;
        RECT 14.85 78.15 15.35 80 ;
        RECT 14.075 78.15 14.575 80 ;
        RECT 13.3 78.15 13.8 80 ;
        RECT 12.525 78.15 13.025 80 ;
        RECT 11.75 78.15 12.25 80 ;
      LAYER C1 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER JA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER QB ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER QA ;
        RECT 12.05 77.975 15.05 80 ;
    END
  END VRES0_B
  PIN VRES3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 72.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.105 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 47.75 78.15 48.25 80 ;
        RECT 46.975 78.15 47.475 80 ;
        RECT 46.2 78.15 46.7 80 ;
        RECT 45.425 78.15 45.925 80 ;
        RECT 44.65 78.15 45.15 80 ;
      LAYER M2 ;
        RECT 47.75 78.15 48.25 80 ;
        RECT 46.975 78.15 47.475 80 ;
        RECT 46.2 78.15 46.7 80 ;
        RECT 45.425 78.15 45.925 80 ;
        RECT 44.65 78.15 45.15 80 ;
      LAYER C1 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER JA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER QB ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER QA ;
        RECT 44.95 77.975 47.95 80 ;
    END
  END VRES3_B
  PIN VESD1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 24.25 78.15 24.75 80 ;
        RECT 23.475 78.15 23.975 80 ;
        RECT 22.7 78.15 23.2 80 ;
        RECT 21.925 78.15 22.425 80 ;
        RECT 21.15 78.15 21.65 80 ;
      LAYER M2 ;
        RECT 24.25 78.15 24.75 80 ;
        RECT 23.475 78.15 23.975 80 ;
        RECT 22.7 78.15 23.2 80 ;
        RECT 21.925 78.15 22.425 80 ;
        RECT 21.15 78.15 21.65 80 ;
      LAYER C1 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER JA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER QB ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER QA ;
        RECT 21.45 77.975 24.45 80 ;
    END
  END VESD1_B
  PIN VRES2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 75.6725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 43.05 78.15 43.55 80 ;
        RECT 42.275 78.15 42.775 80 ;
        RECT 41.5 78.15 42 80 ;
        RECT 40.725 78.15 41.225 80 ;
        RECT 39.95 78.15 40.45 80 ;
      LAYER M2 ;
        RECT 43.05 78.15 43.55 80 ;
        RECT 42.275 78.15 42.775 80 ;
        RECT 41.5 78.15 42 80 ;
        RECT 40.725 78.15 41.225 80 ;
        RECT 39.95 78.15 40.45 80 ;
      LAYER C1 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER JA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER QB ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER QA ;
        RECT 40.25 77.975 43.25 80 ;
    END
  END VRES2_B
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VESD0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 62.855 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 10.15 78.15 10.65 80 ;
        RECT 9.375 78.15 9.875 80 ;
        RECT 8.6 78.15 9.1 80 ;
        RECT 7.825 78.15 8.325 80 ;
        RECT 7.05 78.15 7.55 80 ;
      LAYER M2 ;
        RECT 10.15 78.15 10.65 80 ;
        RECT 9.375 78.15 9.875 80 ;
        RECT 8.6 78.15 9.1 80 ;
        RECT 7.825 78.15 8.325 80 ;
        RECT 7.05 78.15 7.55 80 ;
      LAYER C1 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER JA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER QB ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER QA ;
        RECT 7.35 77.975 10.35 80 ;
    END
  END VESD0_B
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 116.6975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 493.9475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 396.54 LAYER JA ;
    ANTENNAPARTIALMETALAREA 626.15 LAYER QA ;
    ANTENNAPARTIALMETALAREA 396.54 LAYER QB ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 54.72 LAYER JV ;
    ANTENNAPARTIALCUTAREA 54.72 LAYER JW ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A2 ;
    ANTENNADIFFAREA 150.1 LAYER C5 ;
    ANTENNADIFFAREA 150.1 LAYER C4 ;
    ANTENNADIFFAREA 150.1 LAYER JA ;
    ANTENNADIFFAREA 150.1 LAYER QA ;
    ANTENNADIFFAREA 150.1 LAYER QB ;
    ANTENNADIFFAREA 150.1 LAYER C3 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 24 58 28.8 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN VESD2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 38.35 78.15 38.85 80 ;
        RECT 37.575 78.15 38.075 80 ;
        RECT 36.8 78.15 37.3 80 ;
        RECT 36.025 78.15 36.525 80 ;
        RECT 35.25 78.15 35.75 80 ;
      LAYER M2 ;
        RECT 38.35 78.15 38.85 80 ;
        RECT 37.575 78.15 38.075 80 ;
        RECT 36.8 78.15 37.3 80 ;
        RECT 36.025 78.15 36.525 80 ;
        RECT 35.25 78.15 35.75 80 ;
      LAYER C1 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER JA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER QB ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER QA ;
        RECT 35.55 77.975 38.55 80 ;
    END
  END VESD2_B
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_ANACORE_V

MACRO RIIO_EG1D80V_ANAIO_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ANAIO_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VESD3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 63.22955 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 62.855 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 52.45 78.15 52.95 80 ;
        RECT 51.675 78.15 52.175 80 ;
        RECT 50.9 78.15 51.4 80 ;
        RECT 50.125 78.15 50.625 80 ;
        RECT 49.35 78.15 49.85 80 ;
      LAYER M2 ;
        RECT 52.45 78.15 52.95 80 ;
        RECT 51.675 78.15 52.175 80 ;
        RECT 50.9 78.15 51.4 80 ;
        RECT 50.125 78.15 50.625 80 ;
        RECT 49.35 78.15 49.85 80 ;
      LAYER C1 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER JA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER QB ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER QA ;
        RECT 49.65 77.975 52.65 80 ;
    END
  END VESD3_B
  PIN VRES1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 75.6725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 19.55 78.15 20.05 80 ;
        RECT 18.775 78.15 19.275 80 ;
        RECT 18 78.15 18.5 80 ;
        RECT 17.225 78.15 17.725 80 ;
        RECT 16.45 78.15 16.95 80 ;
      LAYER M2 ;
        RECT 19.55 78.15 20.05 80 ;
        RECT 18.775 78.15 19.275 80 ;
        RECT 18 78.15 18.5 80 ;
        RECT 17.225 78.15 17.725 80 ;
        RECT 16.45 78.15 16.95 80 ;
      LAYER C1 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER JA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER QB ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER QA ;
        RECT 16.75 77.975 19.75 80 ;
    END
  END VRES1_B
  PIN VRES0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 72.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 16.735 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.105 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 14.85 78.15 15.35 80 ;
        RECT 14.075 78.15 14.575 80 ;
        RECT 13.3 78.15 13.8 80 ;
        RECT 12.525 78.15 13.025 80 ;
        RECT 11.75 78.15 12.25 80 ;
      LAYER M2 ;
        RECT 14.85 78.15 15.35 80 ;
        RECT 14.075 78.15 14.575 80 ;
        RECT 13.3 78.15 13.8 80 ;
        RECT 12.525 78.15 13.025 80 ;
        RECT 11.75 78.15 12.25 80 ;
      LAYER C1 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER JA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER QB ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER QA ;
        RECT 12.05 77.975 15.05 80 ;
    END
  END VRES0_B
  PIN VRES3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 72.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 10.075 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.105 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 47.75 78.15 48.25 80 ;
        RECT 46.975 78.15 47.475 80 ;
        RECT 46.2 78.15 46.7 80 ;
        RECT 45.425 78.15 45.925 80 ;
        RECT 44.65 78.15 45.15 80 ;
      LAYER M2 ;
        RECT 47.75 78.15 48.25 80 ;
        RECT 46.975 78.15 47.475 80 ;
        RECT 46.2 78.15 46.7 80 ;
        RECT 45.425 78.15 45.925 80 ;
        RECT 44.65 78.15 45.15 80 ;
      LAYER C1 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER JA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER QB ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER QA ;
        RECT 44.95 77.975 47.95 80 ;
    END
  END VRES3_B
  PIN VESD1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 24.25 78.15 24.75 80 ;
        RECT 23.475 78.15 23.975 80 ;
        RECT 22.7 78.15 23.2 80 ;
        RECT 21.925 78.15 22.425 80 ;
        RECT 21.15 78.15 21.65 80 ;
      LAYER M2 ;
        RECT 24.25 78.15 24.75 80 ;
        RECT 23.475 78.15 23.975 80 ;
        RECT 22.7 78.15 23.2 80 ;
        RECT 21.925 78.15 22.425 80 ;
        RECT 21.15 78.15 21.65 80 ;
      LAYER C1 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER JA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER QB ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER QA ;
        RECT 21.45 77.975 24.45 80 ;
    END
  END VESD1_B
  PIN VRES2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 75.6725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 43.05 78.15 43.55 80 ;
        RECT 42.275 78.15 42.775 80 ;
        RECT 41.5 78.15 42 80 ;
        RECT 40.725 78.15 41.225 80 ;
        RECT 39.95 78.15 40.45 80 ;
      LAYER M2 ;
        RECT 43.05 78.15 43.55 80 ;
        RECT 42.275 78.15 42.775 80 ;
        RECT 41.5 78.15 42 80 ;
        RECT 40.725 78.15 41.225 80 ;
        RECT 39.95 78.15 40.45 80 ;
      LAYER C1 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER JA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER QB ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER QA ;
        RECT 40.25 77.975 43.25 80 ;
    END
  END VRES2_B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VESD0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 62.855 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 10.15 78.15 10.65 80 ;
        RECT 9.375 78.15 9.875 80 ;
        RECT 8.6 78.15 9.1 80 ;
        RECT 7.825 78.15 8.325 80 ;
        RECT 7.05 78.15 7.55 80 ;
      LAYER M2 ;
        RECT 10.15 78.15 10.65 80 ;
        RECT 9.375 78.15 9.875 80 ;
        RECT 8.6 78.15 9.1 80 ;
        RECT 7.825 78.15 8.325 80 ;
        RECT 7.05 78.15 7.55 80 ;
      LAYER C1 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER JA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER QB ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER QA ;
        RECT 7.35 77.975 10.35 80 ;
    END
  END VESD0_B
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 116.65125 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 493.90125 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 396.54 LAYER JA ;
    ANTENNAPARTIALMETALAREA 626.15 LAYER QA ;
    ANTENNAPARTIALMETALAREA 396.54 LAYER QB ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 54.72 LAYER JV ;
    ANTENNAPARTIALCUTAREA 54.72 LAYER JW ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A2 ;
    ANTENNADIFFAREA 163.4 LAYER C5 ;
    ANTENNADIFFAREA 163.4 LAYER C4 ;
    ANTENNADIFFAREA 163.4 LAYER JA ;
    ANTENNADIFFAREA 163.4 LAYER QA ;
    ANTENNADIFFAREA 163.4 LAYER QB ;
    ANTENNADIFFAREA 163.4 LAYER C3 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.875 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.875 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER JA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 24 58 28.8 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN VESD2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 38.35 78.15 38.85 80 ;
        RECT 37.575 78.15 38.075 80 ;
        RECT 36.8 78.15 37.3 80 ;
        RECT 36.025 78.15 36.525 80 ;
        RECT 35.25 78.15 35.75 80 ;
      LAYER M2 ;
        RECT 38.35 78.15 38.85 80 ;
        RECT 37.575 78.15 38.075 80 ;
        RECT 36.8 78.15 37.3 80 ;
        RECT 36.025 78.15 36.525 80 ;
        RECT 35.25 78.15 35.75 80 ;
      LAYER C1 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER JA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER QB ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER QA ;
        RECT 35.55 77.975 38.55 80 ;
    END
  END VESD2_B
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_ANAIO_V

MACRO RIIO_EG1D80V_CUTB2B_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTB2B_V 0 0 ;
  SIZE 16 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_r VSSIO_R!" ;
    PORT
      LAYER QB ;
        RECT 8.875 42.6 16 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 8.875 17.8 16 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 8.875 5.4 16 10.2 ;
    END
  END VSSIO_R
  PIN VSS_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_r VSS_R!" ;
    PORT
      LAYER QB ;
        RECT 8.875 67.4 16 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 8.875 48.8 16 53.6 ;
    END
  END VSS_R
  PIN VSSIO_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_l VSSIO_L!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 7.125 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 7.125 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 7.125 10.2 ;
    END
  END VSSIO_L
  PIN VSS_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_l VSS_L!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 7.125 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 7.125 53.6 ;
    END
  END VSS_L
  OBS
    LAYER CA ;
      RECT 0 0 16 80 ;
    LAYER M1 ;
      RECT 0 0 16 80 ;
    LAYER V1 ;
      RECT 0 0 16 80 ;
    LAYER M2 ;
      RECT 0 0 16 80 ;
    LAYER A1 ;
      RECT 0 0 16 80 ;
    LAYER C2 ;
      RECT 0 0 16 80 ;
    LAYER CB ;
      RECT 0 0 16 80 ;
    LAYER JV ;
      RECT 0 0 16 80 ;
    LAYER YS ;
      RECT 0 0 16 80 ;
    LAYER JW ;
      RECT 0 0 16 80 ;
    LAYER QB ;
      RECT 0 0 16 80 ;
    LAYER QA ;
      RECT 0 0 16 80 ;
    LAYER JA ;
      RECT 0 0 16 80 ;
    LAYER AY ;
      RECT 0 0 16 80 ;
    LAYER C1 ;
      RECT 0 0 16 80 ;
    LAYER C5 ;
      RECT 0 0 16 80 ;
    LAYER C4 ;
      RECT 0 0 16 80 ;
    LAYER C3 ;
      RECT 0 0 16 80 ;
    LAYER A4 ;
      RECT 0 0 16 80 ;
    LAYER A3 ;
      RECT 0 0 16 80 ;
    LAYER A2 ;
      RECT 0 0 16 80 ;
  END
END RIIO_EG1D80V_CUTB2B_V

MACRO RIIO_EG1D80V_CUTBIAS_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTBIAS_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 4 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 4 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 4 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 4 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 4 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 4 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 4 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 4 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 4 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 4 53.6 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTBIAS_V

MACRO RIIO_EG1D80V_CUTCOREB2B_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCOREB2B_V 0 0 ;
  SIZE 16 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 16 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 16 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 16 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 16 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 16 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 16 10.2 ;
    END
  END VSSIO
  PIN VSS_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_l VSS_L!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 7.125 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 7.125 53.6 ;
    END
  END VSS_L
  PIN VSS_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_r VSS_R!" ;
    PORT
      LAYER QB ;
        RECT 8.875 67.4 16 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 8.875 48.8 16 53.6 ;
    END
  END VSS_R
  OBS
    LAYER CA ;
      RECT 0 0 16 80 ;
    LAYER M1 ;
      RECT 0 0 16 80 ;
    LAYER V1 ;
      RECT 0 0 16 80 ;
    LAYER M2 ;
      RECT 0 0 16 80 ;
    LAYER A1 ;
      RECT 0 0 16 80 ;
    LAYER C2 ;
      RECT 0 0 16 80 ;
    LAYER CB ;
      RECT 0 0 16 80 ;
    LAYER JV ;
      RECT 0 0 16 80 ;
    LAYER YS ;
      RECT 0 0 16 80 ;
    LAYER JW ;
      RECT 0 0 16 80 ;
    LAYER QB ;
      RECT 0 0 16 80 ;
    LAYER QA ;
      RECT 0 0 16 80 ;
    LAYER JA ;
      RECT 0 0 16 80 ;
    LAYER AY ;
      RECT 0 0 16 80 ;
    LAYER C1 ;
      RECT 0 0 16 80 ;
    LAYER C5 ;
      RECT 0 0 16 80 ;
    LAYER C4 ;
      RECT 0 0 16 80 ;
    LAYER C3 ;
      RECT 0 0 16 80 ;
    LAYER A4 ;
      RECT 0 0 16 80 ;
    LAYER A3 ;
      RECT 0 0 16 80 ;
    LAYER A2 ;
      RECT 0 0 16 80 ;
  END
END RIIO_EG1D80V_CUTCOREB2B_V

MACRO RIIO_EG1D80V_CUTCOREPWR_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCOREPWR_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 4 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 4 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 4 10.2 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 4 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 4 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 4 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 4 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 4 16.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTCOREPWR_V

MACRO RIIO_EG1D80V_CUTCORE_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCORE_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 4 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 4 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 4 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 4 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 4 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 4 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTCORE_V

MACRO RIIO_EG1D80V_CUTIOB2B_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIOB2B_V 0 0 ;
  SIZE 16 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_l VSSIO_L!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 7.125 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 7.125 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 7.125 10.2 ;
    END
  END VSSIO_L
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 16 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 16 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 16 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 16 53.6 ;
    END
  END VSS
  PIN VSSIO_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_r VSSIO_R!" ;
    PORT
      LAYER QB ;
        RECT 8.875 42.6 16 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 8.875 17.8 16 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 8.875 5.4 16 10.2 ;
    END
  END VSSIO_R
  OBS
    LAYER CA ;
      RECT 0 0 16 80 ;
    LAYER M1 ;
      RECT 0 0 16 80 ;
    LAYER V1 ;
      RECT 0 0 16 80 ;
    LAYER M2 ;
      RECT 0 0 16 80 ;
    LAYER A1 ;
      RECT 0 0 16 80 ;
    LAYER C2 ;
      RECT 0 0 16 80 ;
    LAYER CB ;
      RECT 0 0 16 80 ;
    LAYER JV ;
      RECT 0 0 16 80 ;
    LAYER YS ;
      RECT 0 0 16 80 ;
    LAYER JW ;
      RECT 0 0 16 80 ;
    LAYER QB ;
      RECT 0 0 16 80 ;
    LAYER QA ;
      RECT 0 0 16 80 ;
    LAYER JA ;
      RECT 0 0 16 80 ;
    LAYER AY ;
      RECT 0 0 16 80 ;
    LAYER C1 ;
      RECT 0 0 16 80 ;
    LAYER C5 ;
      RECT 0 0 16 80 ;
    LAYER C4 ;
      RECT 0 0 16 80 ;
    LAYER C3 ;
      RECT 0 0 16 80 ;
    LAYER A4 ;
      RECT 0 0 16 80 ;
    LAYER A3 ;
      RECT 0 0 16 80 ;
    LAYER A2 ;
      RECT 0 0 16 80 ;
  END
END RIIO_EG1D80V_CUTIOB2B_V

MACRO RIIO_EG1D80V_CUTIOPWR_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIOPWR_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 4 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 4 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 4 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 4 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 4 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 4 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 4 53.6 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTIOPWR_V

MACRO RIIO_EG1D80V_CUTIO_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIO_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 4 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 4 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 4 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 4 53.6 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTIO_V

MACRO RIIO_EG1D80V_CUTPWR_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTPWR_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 4 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 4 53.6 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 4 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 4 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 4 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTPWR_V

MACRO RIIO_EG1D80V_CUT_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUT_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUT_V

MACRO RIIO_EG1D80V_FILL16B2B_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL16B2B_V 0 0 ;
  SIZE 16 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 16 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 16 53.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 16 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 16 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 16 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 16 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 16 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 16 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 16 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 16 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 16 80 ;
    LAYER M1 ;
      RECT 0 0 16 80 ;
    LAYER V1 ;
      RECT 0 0 16 80 ;
    LAYER M2 ;
      RECT 0 0 16 80 ;
    LAYER A1 ;
      RECT 0 0 16 80 ;
    LAYER C2 ;
      RECT 0 0 16 80 ;
    LAYER CB ;
      RECT 0 0 16 80 ;
    LAYER JV ;
      RECT 0 0 16 80 ;
    LAYER YS ;
      RECT 0 0 16 80 ;
    LAYER JW ;
      RECT 0 0 16 80 ;
    LAYER QB ;
      RECT 0 0 16 80 ;
    LAYER QA ;
      RECT 0 0 16 80 ;
    LAYER JA ;
      RECT 0 0 16 80 ;
    LAYER AY ;
      RECT 0 0 16 80 ;
    LAYER C1 ;
      RECT 0 0 16 80 ;
    LAYER C5 ;
      RECT 0 0 16 80 ;
    LAYER C4 ;
      RECT 0 0 16 80 ;
    LAYER C3 ;
      RECT 0 0 16 80 ;
    LAYER A4 ;
      RECT 0 0 16 80 ;
    LAYER A3 ;
      RECT 0 0 16 80 ;
    LAYER A2 ;
      RECT 0 0 16 80 ;
  END
END RIIO_EG1D80V_FILL16B2B_V

MACRO RIIO_EG1D80V_FILL16_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL16_V 0 0 ;
  SIZE 16 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 16 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 16 53.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 16 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 16 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 16 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 16 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 16 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 16 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 16 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 16 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 16 80 ;
    LAYER M1 ;
      RECT 0 0 16 80 ;
    LAYER V1 ;
      RECT 0 0 16 80 ;
    LAYER M2 ;
      RECT 0 0 16 80 ;
    LAYER A1 ;
      RECT 0 0 16 80 ;
    LAYER C2 ;
      RECT 0 0 16 80 ;
    LAYER CB ;
      RECT 0 0 16 80 ;
    LAYER JV ;
      RECT 0 0 16 80 ;
    LAYER YS ;
      RECT 0 0 16 80 ;
    LAYER JW ;
      RECT 0 0 16 80 ;
    LAYER QB ;
      RECT 0 0 16 80 ;
    LAYER QA ;
      RECT 0 0 16 80 ;
    LAYER JA ;
      RECT 0 0 16 80 ;
    LAYER AY ;
      RECT 0 0 16 80 ;
    LAYER C1 ;
      RECT 0 0 16 80 ;
    LAYER C5 ;
      RECT 0 0 16 80 ;
    LAYER C4 ;
      RECT 0 0 16 80 ;
    LAYER C3 ;
      RECT 0 0 16 80 ;
    LAYER A4 ;
      RECT 0 0 16 80 ;
    LAYER A3 ;
      RECT 0 0 16 80 ;
    LAYER A2 ;
      RECT 0 0 16 80 ;
  END
END RIIO_EG1D80V_FILL16_V

MACRO RIIO_EG1D80V_FILL1_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL1_V 0 0 ;
  SIZE 1 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 1 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 1 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 1 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 1 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 1 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 1 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 1 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 1 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 1 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 1 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 1 80 ;
    LAYER M1 ;
      RECT 0 0 1 80 ;
    LAYER V1 ;
      RECT 0 0 1 80 ;
    LAYER M2 ;
      RECT 0 0 1 80 ;
    LAYER A1 ;
      RECT 0 0 1 80 ;
    LAYER C2 ;
      RECT 0 0 1 80 ;
    LAYER CB ;
      RECT 0 0 1 80 ;
    LAYER JV ;
      RECT 0 0 1 80 ;
    LAYER YS ;
      RECT 0 0 1 80 ;
    LAYER JW ;
      RECT 0 0 1 80 ;
    LAYER QB ;
      RECT 0 0 1 80 ;
    LAYER QA ;
      RECT 0 0 1 80 ;
    LAYER JA ;
      RECT 0 0 1 80 ;
    LAYER AY ;
      RECT 0 0 1 80 ;
    LAYER C1 ;
      RECT 0 0 1 80 ;
    LAYER C5 ;
      RECT 0 0 1 80 ;
    LAYER C4 ;
      RECT 0 0 1 80 ;
    LAYER C3 ;
      RECT 0 0 1 80 ;
    LAYER A4 ;
      RECT 0 0 1 80 ;
    LAYER A3 ;
      RECT 0 0 1 80 ;
    LAYER A2 ;
      RECT 0 0 1 80 ;
  END
END RIIO_EG1D80V_FILL1_V

MACRO RIIO_EG1D80V_FILL2_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL2_V 0 0 ;
  SIZE 2 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 2 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 2 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 2 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 2 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 2 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 2 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 2 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 2 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 2 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 2 16.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 2 80 ;
    LAYER M1 ;
      RECT 0 0 2 80 ;
    LAYER V1 ;
      RECT 0 0 2 80 ;
    LAYER M2 ;
      RECT 0 0 2 80 ;
    LAYER A1 ;
      RECT 0 0 2 80 ;
    LAYER C2 ;
      RECT 0 0 2 80 ;
    LAYER CB ;
      RECT 0 0 2 80 ;
    LAYER JV ;
      RECT 0 0 2 80 ;
    LAYER YS ;
      RECT 0 0 2 80 ;
    LAYER JW ;
      RECT 0 0 2 80 ;
    LAYER QB ;
      RECT 0 0 2 80 ;
    LAYER QA ;
      RECT 0 0 2 80 ;
    LAYER JA ;
      RECT 0 0 2 80 ;
    LAYER AY ;
      RECT 0 0 2 80 ;
    LAYER C1 ;
      RECT 0 0 2 80 ;
    LAYER C5 ;
      RECT 0 0 2 80 ;
    LAYER C4 ;
      RECT 0 0 2 80 ;
    LAYER C3 ;
      RECT 0 0 2 80 ;
    LAYER A4 ;
      RECT 0 0 2 80 ;
    LAYER A3 ;
      RECT 0 0 2 80 ;
    LAYER A2 ;
      RECT 0 0 2 80 ;
  END
END RIIO_EG1D80V_FILL2_V

MACRO RIIO_EG1D80V_FILL32_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL32_V 0 0 ;
  SIZE 32 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 32 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 32 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 32 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 32 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 32 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 32 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 32 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 32 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 32 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 32 53.6 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 32 80 ;
    LAYER M1 ;
      RECT 0 0 32 80 ;
    LAYER V1 ;
      RECT 0 0 32 80 ;
    LAYER M2 ;
      RECT 0 0 32 80 ;
    LAYER A1 ;
      RECT 0 0 32 80 ;
    LAYER C2 ;
      RECT 0 0 32 80 ;
    LAYER CB ;
      RECT 0 0 32 80 ;
    LAYER JV ;
      RECT 0 0 32 80 ;
    LAYER YS ;
      RECT 0 0 32 80 ;
    LAYER JW ;
      RECT 0 0 32 80 ;
    LAYER QB ;
      RECT 0 0 32 80 ;
    LAYER QA ;
      RECT 0 0 32 80 ;
    LAYER JA ;
      RECT 0 0 32 80 ;
    LAYER AY ;
      RECT 0 0 32 80 ;
    LAYER C1 ;
      RECT 0 0 32 80 ;
    LAYER C5 ;
      RECT 0 0 32 80 ;
    LAYER C4 ;
      RECT 0 0 32 80 ;
    LAYER C3 ;
      RECT 0 0 32 80 ;
    LAYER A4 ;
      RECT 0 0 32 80 ;
    LAYER A3 ;
      RECT 0 0 32 80 ;
    LAYER A2 ;
      RECT 0 0 32 80 ;
  END
END RIIO_EG1D80V_FILL32_V

MACRO RIIO_EG1D80V_FILL4_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL4_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 4 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 4 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 4 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 4 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 4 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 4 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 4 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 4 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 4 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 4 53.6 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_FILL4_V

MACRO RIIO_EG1D80V_FILL8_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL8_V 0 0 ;
  SIZE 8 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 8 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 8 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 8 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 8 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 8 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 8 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 8 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 8 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 8 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 8 53.6 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 8 80 ;
    LAYER M1 ;
      RECT 0 0 8 80 ;
    LAYER V1 ;
      RECT 0 0 8 80 ;
    LAYER M2 ;
      RECT 0 0 8 80 ;
    LAYER A1 ;
      RECT 0 0 8 80 ;
    LAYER C2 ;
      RECT 0 0 8 80 ;
    LAYER CB ;
      RECT 0 0 8 80 ;
    LAYER JV ;
      RECT 0 0 8 80 ;
    LAYER YS ;
      RECT 0 0 8 80 ;
    LAYER JW ;
      RECT 0 0 8 80 ;
    LAYER QB ;
      RECT 0 0 8 80 ;
    LAYER QA ;
      RECT 0 0 8 80 ;
    LAYER JA ;
      RECT 0 0 8 80 ;
    LAYER AY ;
      RECT 0 0 8 80 ;
    LAYER C1 ;
      RECT 0 0 8 80 ;
    LAYER C5 ;
      RECT 0 0 8 80 ;
    LAYER C4 ;
      RECT 0 0 8 80 ;
    LAYER C3 ;
      RECT 0 0 8 80 ;
    LAYER A4 ;
      RECT 0 0 8 80 ;
    LAYER A3 ;
      RECT 0 0 8 80 ;
    LAYER A2 ;
      RECT 0 0 8 80 ;
  END
END RIIO_EG1D80V_FILL8_V

MACRO RIIO_EG1D80V_POR_IO_V1D0_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_POR_IO_V1D0_V 0 0 ;
  SIZE 8 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER C2 ;
        RECT 0 37.075 8 39.575 ;
    END
    PORT
      LAYER QB ;
        RECT 0 42.6 8 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 8 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 8 10.2 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER C2 ;
        RECT 0 74.575 8 77.075 ;
    END
    PORT
      LAYER QB ;
        RECT 0 67.4 8 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 8 53.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER C2 ;
        RECT 0 70.825 8 73.325 ;
    END
    PORT
      LAYER QB ;
        RECT 0 61.2 8 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 8 59.8 ;
    END
  END VDD
  PIN VDDIO_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio_por VDDIO_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 1.25 33.325 1.75 80 ;
    END
  END VDDIO_POR
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 8 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 8 35 ;
      LAYER C2 ;
        RECT 0 33.325 8 35.825 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 8 16.4 ;
    END
  END VDDIO
  PIN VSSIO_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_por VSSIO_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 2.25 33.325 2.75 80 ;
    END
  END VSSIO_POR
  PIN POR_N_CORE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.5875 LAYER C1 ;
    ANTENNADIFFAREA 0.3135 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.25 79.5 6.75 80 ;
    END
  END POR_N_CORE_O
  PIN VDD_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd_por VDD_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 5.25 70.825 5.75 80 ;
    END
  END VDD_POR
  PIN VSS_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_por VSS_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 4.25 70.825 4.75 80 ;
    END
  END VSS_POR
  OBS
    LAYER CA ;
      RECT 0 0 8 80 ;
    LAYER M1 ;
      RECT 0 0 8 80 ;
    LAYER V1 ;
      RECT 0 0 8 80 ;
    LAYER M2 ;
      RECT 0 0 8 80 ;
    LAYER A1 ;
      RECT 0 0 8 80 ;
    LAYER C2 ;
      RECT 0 0 8 80 ;
    LAYER CB ;
      RECT 0 0 8 80 ;
    LAYER JV ;
      RECT 0 0 8 80 ;
    LAYER YS ;
      RECT 0 0 8 80 ;
    LAYER JW ;
      RECT 0 0 8 80 ;
    LAYER QB ;
      RECT 0 0 8 80 ;
    LAYER QA ;
      RECT 0 0 8 80 ;
    LAYER JA ;
      RECT 0 0 8 80 ;
    LAYER AY ;
      RECT 0 0 8 80 ;
    LAYER C1 ;
      RECT 0 0 8 80 ;
    LAYER C5 ;
      RECT 0 0 8 80 ;
    LAYER C4 ;
      RECT 0 0 8 80 ;
    LAYER C3 ;
      RECT 0 0 8 80 ;
    LAYER A4 ;
      RECT 0 0 8 80 ;
    LAYER A3 ;
      RECT 0 0 8 80 ;
    LAYER A2 ;
      RECT 0 0 8 80 ;
  END
END RIIO_EG1D80V_POR_IO_V1D0_V

MACRO RIIO_EG1D80V_RAILSHORT_GND_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_GND_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 4 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 4 53.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 42.6 4 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 4 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 4 10.2 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 4 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 4 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 4 16.4 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 4 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 4 59.8 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_RAILSHORT_GND_V

MACRO RIIO_EG1D80V_RAILSHORT_PG_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_PG_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 4 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 4 59.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 36.4 4 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 4 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 4 16.4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 4 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 4 53.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 42.6 4 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 4 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 4 10.2 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_RAILSHORT_PG_V

MACRO RIIO_EG1D80V_RAILSHORT_PWR_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_PWR_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 4 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 4 59.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 36.4 4 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 4 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 4 16.4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 4 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 4 53.6 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 4 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 4 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 4 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER JV ;
      RECT 0 0 4 80 ;
    LAYER YS ;
      RECT 0 0 4 80 ;
    LAYER JW ;
      RECT 0 0 4 80 ;
    LAYER QB ;
      RECT 0 0 4 80 ;
    LAYER QA ;
      RECT 0 0 4 80 ;
    LAYER JA ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_RAILSHORT_PWR_V

MACRO RIIO_EG1D80V_VDD04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
    END
    PORT
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
    END
    PORT
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
    END
    PORT
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDD04_V

MACRO RIIO_EG1D80V_VDDIOX_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDIOX_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSSIOX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssiox VSSIOX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
        RECT 9.837 79.19 12.662 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 47.337 79.19 50.162 80 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
  END VSSIOX
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDDIOX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddiox VDDIOX!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VDDIOX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDIOX_V

MACRO RIIO_EG1D80V_VDDIO_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDIO_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDIO_V

MACRO RIIO_EG1D80V_VDDQ04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSQ
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VDDQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDQ04_V

MACRO RIIO_EG1D80V_VDDQ_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VDDQ
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDQ_HVT_V

MACRO RIIO_EG1D80V_VDDQ_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VDDQ
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDQ_RVT_V

MACRO RIIO_EG1D80V_VDDX04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.25 78.15 8.75 80 ;
        RECT 2.5 78.15 5 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.25 78.15 8.75 80 ;
        RECT 2.5 78.15 5 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
        RECT 9.837 79.19 12.662 80 ;
        RECT 6.087 79.19 8.912 80 ;
        RECT 2.337 79.19 5.162 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.412 79.19 8.912 80 ;
        RECT 7.637 79.19 8.137 80 ;
        RECT 6.862 79.19 7.362 80 ;
        RECT 6.087 79.19 6.587 80 ;
        RECT 4.662 79.19 5.162 80 ;
        RECT 3.887 79.19 4.387 80 ;
        RECT 3.112 79.19 3.612 80 ;
        RECT 2.337 79.19 2.837 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.412 79.19 8.912 80 ;
        RECT 7.637 79.19 8.137 80 ;
        RECT 6.862 79.19 7.362 80 ;
        RECT 6.087 79.19 6.587 80 ;
        RECT 4.662 79.19 5.162 80 ;
        RECT 3.887 79.19 4.387 80 ;
        RECT 3.112 79.19 3.612 80 ;
        RECT 2.337 79.19 2.837 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 55 78.15 57.5 80 ;
        RECT 51.25 78.15 53.75 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 55 78.15 57.5 80 ;
        RECT 51.25 78.15 53.75 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 54.837 79.19 57.662 80 ;
        RECT 51.087 79.19 53.912 80 ;
        RECT 47.337 79.19 50.162 80 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M1 ;
        RECT 57.162 79.19 57.662 80 ;
        RECT 56.387 79.19 56.887 80 ;
        RECT 55.612 79.19 56.112 80 ;
        RECT 54.837 79.19 55.337 80 ;
        RECT 53.412 79.19 53.912 80 ;
        RECT 52.637 79.19 53.137 80 ;
        RECT 51.862 79.19 52.362 80 ;
        RECT 51.087 79.19 51.587 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M2 ;
        RECT 57.162 79.19 57.662 80 ;
        RECT 56.387 79.19 56.887 80 ;
        RECT 55.612 79.19 56.112 80 ;
        RECT 54.837 79.19 55.337 80 ;
        RECT 53.412 79.19 53.912 80 ;
        RECT 52.637 79.19 53.137 80 ;
        RECT 51.862 79.19 52.362 80 ;
        RECT 51.087 79.19 51.587 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDX04_V

MACRO RIIO_EG1D80V_VDDX_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.25 78.15 8.75 80 ;
        RECT 2.5 78.15 5 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.25 78.15 8.75 80 ;
        RECT 2.5 78.15 5 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
        RECT 9.837 79.19 12.662 80 ;
        RECT 6.087 79.19 8.912 80 ;
        RECT 2.337 79.19 5.162 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.412 79.19 8.912 80 ;
        RECT 7.637 79.19 8.137 80 ;
        RECT 6.862 79.19 7.362 80 ;
        RECT 6.087 79.19 6.587 80 ;
        RECT 4.662 79.19 5.162 80 ;
        RECT 3.887 79.19 4.387 80 ;
        RECT 3.112 79.19 3.612 80 ;
        RECT 2.337 79.19 2.837 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.412 79.19 8.912 80 ;
        RECT 7.637 79.19 8.137 80 ;
        RECT 6.862 79.19 7.362 80 ;
        RECT 6.087 79.19 6.587 80 ;
        RECT 4.662 79.19 5.162 80 ;
        RECT 3.887 79.19 4.387 80 ;
        RECT 3.112 79.19 3.612 80 ;
        RECT 2.337 79.19 2.837 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 55 78.15 57.5 80 ;
        RECT 51.25 78.15 53.75 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 55 78.15 57.5 80 ;
        RECT 51.25 78.15 53.75 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 54.837 79.19 57.662 80 ;
        RECT 51.087 79.19 53.912 80 ;
        RECT 47.337 79.19 50.162 80 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 57.162 79.19 57.662 80 ;
        RECT 56.387 79.19 56.887 80 ;
        RECT 55.612 79.19 56.112 80 ;
        RECT 54.837 79.19 55.337 80 ;
        RECT 53.412 79.19 53.912 80 ;
        RECT 52.637 79.19 53.137 80 ;
        RECT 51.862 79.19 52.362 80 ;
        RECT 51.087 79.19 51.587 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 57.162 79.19 57.662 80 ;
        RECT 56.387 79.19 56.887 80 ;
        RECT 55.612 79.19 56.112 80 ;
        RECT 54.837 79.19 55.337 80 ;
        RECT 53.412 79.19 53.912 80 ;
        RECT 52.637 79.19 53.137 80 ;
        RECT 51.862 79.19 52.362 80 ;
        RECT 51.087 79.19 51.587 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDX_HVT_V

MACRO RIIO_EG1D80V_VDDX_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.25 78.15 8.75 80 ;
        RECT 2.5 78.15 5 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.25 78.15 8.75 80 ;
        RECT 2.5 78.15 5 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
        RECT 9.837 79.19 12.662 80 ;
        RECT 6.087 79.19 8.912 80 ;
        RECT 2.337 79.19 5.162 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.412 79.19 8.912 80 ;
        RECT 7.637 79.19 8.137 80 ;
        RECT 6.862 79.19 7.362 80 ;
        RECT 6.087 79.19 6.587 80 ;
        RECT 4.662 79.19 5.162 80 ;
        RECT 3.887 79.19 4.387 80 ;
        RECT 3.112 79.19 3.612 80 ;
        RECT 2.337 79.19 2.837 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.412 79.19 8.912 80 ;
        RECT 7.637 79.19 8.137 80 ;
        RECT 6.862 79.19 7.362 80 ;
        RECT 6.087 79.19 6.587 80 ;
        RECT 4.662 79.19 5.162 80 ;
        RECT 3.887 79.19 4.387 80 ;
        RECT 3.112 79.19 3.612 80 ;
        RECT 2.337 79.19 2.837 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 55 78.15 57.5 80 ;
        RECT 51.25 78.15 53.75 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 55 78.15 57.5 80 ;
        RECT 51.25 78.15 53.75 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 54.837 79.19 57.662 80 ;
        RECT 51.087 79.19 53.912 80 ;
        RECT 47.337 79.19 50.162 80 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 57.162 79.19 57.662 80 ;
        RECT 56.387 79.19 56.887 80 ;
        RECT 55.612 79.19 56.112 80 ;
        RECT 54.837 79.19 55.337 80 ;
        RECT 53.412 79.19 53.912 80 ;
        RECT 52.637 79.19 53.137 80 ;
        RECT 51.862 79.19 52.362 80 ;
        RECT 51.087 79.19 51.587 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 57.162 79.19 57.662 80 ;
        RECT 56.387 79.19 56.887 80 ;
        RECT 55.612 79.19 56.112 80 ;
        RECT 54.837 79.19 55.337 80 ;
        RECT 53.412 79.19 53.912 80 ;
        RECT 52.637 79.19 53.137 80 ;
        RECT 51.862 79.19 52.362 80 ;
        RECT 51.087 79.19 51.587 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDX_RVT_V

MACRO RIIO_EG1D80V_VDD_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDD_HVT_V

MACRO RIIO_EG1D80V_VDD_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDD_RVT_V

MACRO RIIO_EG1D80V_VNWINT_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNWINT_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VNWINT_HVT_V

MACRO RIIO_EG1D80V_VNWINT_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNWINT_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VNWINT_RVT_V

MACRO RIIO_EG1D80V_VNW_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNW_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VNW_V

MACRO RIIO_EG1D80V_VPWINT_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPWINT_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VPWINT_HVT_V

MACRO RIIO_EG1D80V_VPWINT_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPWINT_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VPWINT_RVT_V

MACRO RIIO_EG1D80V_VPW_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPW_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VPW_V

MACRO RIIO_EG1D80V_VSS04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSS04_V

MACRO RIIO_EG1D80V_VSSIOX_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSIOX_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSIOX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssiox VSSIOX!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.249 78.15 8.749 80 ;
        RECT 2.498 78.15 4.998 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.249 78.15 8.749 80 ;
        RECT 2.498 78.15 4.998 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
        RECT 9.837 79.19 12.662 80 ;
        RECT 6.086 79.19 8.911 80 ;
        RECT 2.335 79.19 5.16 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.411 79.19 8.911 80 ;
        RECT 7.636 79.19 8.136 80 ;
        RECT 6.861 79.19 7.361 80 ;
        RECT 6.086 79.19 6.586 80 ;
        RECT 4.66 79.19 5.16 80 ;
        RECT 3.885 79.19 4.385 80 ;
        RECT 3.11 79.19 3.61 80 ;
        RECT 2.335 79.19 2.835 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.411 79.19 8.911 80 ;
        RECT 7.636 79.19 8.136 80 ;
        RECT 6.861 79.19 7.361 80 ;
        RECT 6.086 79.19 6.586 80 ;
        RECT 4.66 79.19 5.16 80 ;
        RECT 3.885 79.19 4.385 80 ;
        RECT 3.11 79.19 3.61 80 ;
        RECT 2.335 79.19 2.835 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 54.998 78.15 57.498 80 ;
        RECT 51.249 78.15 53.749 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 54.998 78.15 57.498 80 ;
        RECT 51.249 78.15 53.749 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 54.835 79.19 57.66 80 ;
        RECT 51.086 79.19 53.911 80 ;
        RECT 47.337 79.19 50.162 80 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 57.16 79.19 57.66 80 ;
        RECT 56.385 79.19 56.885 80 ;
        RECT 55.61 79.19 56.11 80 ;
        RECT 54.835 79.19 55.335 80 ;
        RECT 53.411 79.19 53.911 80 ;
        RECT 52.636 79.19 53.136 80 ;
        RECT 51.861 79.19 52.361 80 ;
        RECT 51.086 79.19 51.586 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 57.16 79.19 57.66 80 ;
        RECT 56.385 79.19 56.885 80 ;
        RECT 55.61 79.19 56.11 80 ;
        RECT 54.835 79.19 55.335 80 ;
        RECT 53.411 79.19 53.911 80 ;
        RECT 52.636 79.19 53.136 80 ;
        RECT 51.861 79.19 52.361 80 ;
        RECT 51.086 79.19 51.586 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VSSIOX
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDDIOX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddiox VDDIOX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
    END
  END VDDIOX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSIOX_V

MACRO RIIO_EG1D80V_VSSIO_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSIO_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSIO_V

MACRO RIIO_EG1D80V_VSSQ04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDQ
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VSSQ
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSQ04_V

MACRO RIIO_EG1D80V_VSSQ_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VSSQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSQ_HVT_V

MACRO RIIO_EG1D80V_VSSQ_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VSSQ
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSQ_RVT_V

MACRO RIIO_EG1D80V_VSSX04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.249 78.15 8.749 80 ;
        RECT 2.499 78.15 4.999 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.249 78.15 8.749 80 ;
        RECT 2.499 78.15 4.999 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
        RECT 9.837 79.19 12.662 80 ;
        RECT 6.086 79.19 8.911 80 ;
        RECT 2.336 79.19 5.161 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.411 79.19 8.911 80 ;
        RECT 7.636 79.19 8.136 80 ;
        RECT 6.861 79.19 7.361 80 ;
        RECT 6.086 79.19 6.586 80 ;
        RECT 4.661 79.19 5.161 80 ;
        RECT 3.886 79.19 4.386 80 ;
        RECT 3.111 79.19 3.611 80 ;
        RECT 2.336 79.19 2.836 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.411 79.19 8.911 80 ;
        RECT 7.636 79.19 8.136 80 ;
        RECT 6.861 79.19 7.361 80 ;
        RECT 6.086 79.19 6.586 80 ;
        RECT 4.661 79.19 5.161 80 ;
        RECT 3.886 79.19 4.386 80 ;
        RECT 3.111 79.19 3.611 80 ;
        RECT 2.336 79.19 2.836 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 54.997 78.15 57.497 80 ;
        RECT 51.248 78.15 53.748 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 54.997 78.15 57.497 80 ;
        RECT 51.248 78.15 53.748 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 54.834 79.19 57.659 80 ;
        RECT 51.085 79.19 53.91 80 ;
        RECT 47.337 79.19 50.162 80 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M1 ;
        RECT 57.159 79.19 57.659 80 ;
        RECT 56.384 79.19 56.884 80 ;
        RECT 55.609 79.19 56.109 80 ;
        RECT 54.834 79.19 55.334 80 ;
        RECT 53.41 79.19 53.91 80 ;
        RECT 52.635 79.19 53.135 80 ;
        RECT 51.86 79.19 52.36 80 ;
        RECT 51.085 79.19 51.585 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M2 ;
        RECT 57.159 79.19 57.659 80 ;
        RECT 56.384 79.19 56.884 80 ;
        RECT 55.609 79.19 56.109 80 ;
        RECT 54.834 79.19 55.334 80 ;
        RECT 53.41 79.19 53.91 80 ;
        RECT 52.635 79.19 53.135 80 ;
        RECT 51.86 79.19 52.36 80 ;
        RECT 51.085 79.19 51.585 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSX04_V

MACRO RIIO_EG1D80V_VSSX_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.249 78.15 8.749 80 ;
        RECT 2.499 78.15 4.999 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.249 78.15 8.749 80 ;
        RECT 2.499 78.15 4.999 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
        RECT 9.837 79.19 12.662 80 ;
        RECT 6.086 79.19 8.911 80 ;
        RECT 2.336 79.19 5.161 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.411 79.19 8.911 80 ;
        RECT 7.636 79.19 8.136 80 ;
        RECT 6.861 79.19 7.361 80 ;
        RECT 6.086 79.19 6.586 80 ;
        RECT 4.661 79.19 5.161 80 ;
        RECT 3.886 79.19 4.386 80 ;
        RECT 3.111 79.19 3.611 80 ;
        RECT 2.336 79.19 2.836 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.411 79.19 8.911 80 ;
        RECT 7.636 79.19 8.136 80 ;
        RECT 6.861 79.19 7.361 80 ;
        RECT 6.086 79.19 6.586 80 ;
        RECT 4.661 79.19 5.161 80 ;
        RECT 3.886 79.19 4.386 80 ;
        RECT 3.111 79.19 3.611 80 ;
        RECT 2.336 79.19 2.836 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 54.997 78.15 57.497 80 ;
        RECT 51.248 78.15 53.748 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 54.997 78.15 57.497 80 ;
        RECT 51.248 78.15 53.748 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 54.834 79.19 57.659 80 ;
        RECT 51.085 79.19 53.91 80 ;
        RECT 47.337 79.19 50.162 80 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 57.159 79.19 57.659 80 ;
        RECT 56.384 79.19 56.884 80 ;
        RECT 55.609 79.19 56.109 80 ;
        RECT 54.834 79.19 55.334 80 ;
        RECT 53.41 79.19 53.91 80 ;
        RECT 52.635 79.19 53.135 80 ;
        RECT 51.86 79.19 52.36 80 ;
        RECT 51.085 79.19 51.585 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 57.159 79.19 57.659 80 ;
        RECT 56.384 79.19 56.884 80 ;
        RECT 55.609 79.19 56.109 80 ;
        RECT 54.834 79.19 55.334 80 ;
        RECT 53.41 79.19 53.91 80 ;
        RECT 52.635 79.19 53.135 80 ;
        RECT 51.86 79.19 52.36 80 ;
        RECT 51.085 79.19 51.585 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSX_HVT_V

MACRO RIIO_EG1D80V_VSSX_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.249 78.15 8.749 80 ;
        RECT 2.499 78.15 4.999 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
        RECT 10 78.15 12.5 80 ;
        RECT 6.249 78.15 8.749 80 ;
        RECT 2.499 78.15 4.999 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
        RECT 9.837 79.19 12.662 80 ;
        RECT 6.086 79.19 8.911 80 ;
        RECT 2.336 79.19 5.161 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.411 79.19 8.911 80 ;
        RECT 7.636 79.19 8.136 80 ;
        RECT 6.861 79.19 7.361 80 ;
        RECT 6.086 79.19 6.586 80 ;
        RECT 4.661 79.19 5.161 80 ;
        RECT 3.886 79.19 4.386 80 ;
        RECT 3.111 79.19 3.611 80 ;
        RECT 2.336 79.19 2.836 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
        RECT 8.411 79.19 8.911 80 ;
        RECT 7.636 79.19 8.136 80 ;
        RECT 6.861 79.19 7.361 80 ;
        RECT 6.086 79.19 6.586 80 ;
        RECT 4.661 79.19 5.161 80 ;
        RECT 3.886 79.19 4.386 80 ;
        RECT 3.111 79.19 3.611 80 ;
        RECT 2.336 79.19 2.836 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 54.997 78.15 57.497 80 ;
        RECT 51.248 78.15 53.748 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 54.997 78.15 57.497 80 ;
        RECT 51.248 78.15 53.748 80 ;
        RECT 47.5 78.15 50 80 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 54.834 79.19 57.659 80 ;
        RECT 51.085 79.19 53.91 80 ;
        RECT 47.337 79.19 50.162 80 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 57.159 79.19 57.659 80 ;
        RECT 56.384 79.19 56.884 80 ;
        RECT 55.609 79.19 56.109 80 ;
        RECT 54.834 79.19 55.334 80 ;
        RECT 53.41 79.19 53.91 80 ;
        RECT 52.635 79.19 53.135 80 ;
        RECT 51.86 79.19 52.36 80 ;
        RECT 51.085 79.19 51.585 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 57.159 79.19 57.659 80 ;
        RECT 56.384 79.19 56.884 80 ;
        RECT 55.609 79.19 56.109 80 ;
        RECT 54.834 79.19 55.334 80 ;
        RECT 53.41 79.19 53.91 80 ;
        RECT 52.635 79.19 53.135 80 ;
        RECT 51.86 79.19 52.36 80 ;
        RECT 51.085 79.19 51.585 80 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER QB ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER JA ;
        RECT 27.6 75.2 32.4 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER QB ;
        RECT 27.6 75.2 32.4 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSX_RVT_V

MACRO RIIO_EG1D80V_VSS_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSS_HVT_V

MACRO RIIO_EG1D80V_VSS_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
    END
    PORT
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
    END
    PORT
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
    END
    PORT
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
    END
    PORT
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSS_RVT_V

MACRO RIIO_EG1D80V_VSUP_CORE_GND_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_GND_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSUP
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_CORE_GND_V

MACRO RIIO_EG1D80V_VSUP_CORE_PWR_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_PWR_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSUP
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_CORE_PWR_V

MACRO RIIO_EG1D80V_VSUP_CORE_SIG_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_SIG_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1201.173 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 4.4055 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 514.88 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 1152.81 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 610.4525 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 949.665 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 660.48 LAYER JA ;
    ANTENNAPARTIALMETALAREA 1735.68 LAYER QA ;
    ANTENNAPARTIALMETALAREA 660.48 LAYER QB ;
    ANTENNAPARTIALMETALAREA 4.554 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 18.283584 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 1.792 LAYER AY ;
    ANTENNAPARTIALCUTAREA 16.239168 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 46.27692 LAYER YS ;
    ANTENNAPARTIALCUTAREA 106.56 LAYER JV ;
    ANTENNAPARTIALCUTAREA 106.56 LAYER JW ;
    ANTENNAPARTIALCUTAREA 1.92 LAYER V1 ;
    ANTENNADIFFAREA 150.1 LAYER C3 ;
    ANTENNADIFFAREA 150.1 LAYER C2 ;
    ANTENNADIFFAREA 150.1 LAYER C4 ;
    ANTENNADIFFAREA 150.1 LAYER C5 ;
    ANTENNADIFFAREA 150.1 LAYER JA ;
    ANTENNADIFFAREA 150.1 LAYER QA ;
    ANTENNADIFFAREA 150.1 LAYER QB ;
    ANTENNADIFFAREA 150.1 LAYER C1 ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
        RECT 2.65 79.19 5.65 80 ;
    END
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
        RECT 2 24 58 28.8 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END VSUP
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_CORE_SIG_V

MACRO RIIO_EG1D80V_VSUP_IO_GND_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_GND_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSUP
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_IO_GND_V

MACRO RIIO_EG1D80V_VSUP_IO_PWR_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_PWR_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER QA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER JA ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER QB ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER QA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER JA ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER QA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER JA ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER QB ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER QA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER JA ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER QA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER JA ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER QB ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER QA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER JA ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER QB ;
        RECT 2 24 58 28.8 ;
    END
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSUP
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_IO_PWR_V

MACRO RIIO_EG1D80V_VSUP_IO_SIG_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_SIG_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1543.173 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 4.4055 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 654.255 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 1152.81 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 610.4525 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 949.665 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 660.48 LAYER JA ;
    ANTENNAPARTIALMETALAREA 1735.68 LAYER QA ;
    ANTENNAPARTIALMETALAREA 660.48 LAYER QB ;
    ANTENNAPARTIALMETALAREA 4.554 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 23.58048 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 1.792 LAYER AY ;
    ANTENNAPARTIALCUTAREA 19.220608 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 46.27692 LAYER YS ;
    ANTENNAPARTIALCUTAREA 106.56 LAYER JV ;
    ANTENNAPARTIALCUTAREA 106.56 LAYER JW ;
    ANTENNAPARTIALCUTAREA 1.92 LAYER V1 ;
    ANTENNADIFFAREA 163.4 LAYER C3 ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    ANTENNADIFFAREA 163.4 LAYER C4 ;
    ANTENNADIFFAREA 163.4 LAYER C5 ;
    ANTENNADIFFAREA 163.4 LAYER JA ;
    ANTENNADIFFAREA 163.4 LAYER QA ;
    ANTENNADIFFAREA 163.4 LAYER QB ;
    ANTENNADIFFAREA 163.4 LAYER C1 ;
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER QA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER JA ;
        RECT 53.2 75.2 58 80 ;
        RECT 46.8 75.2 51.6 80 ;
        RECT 40.4 75.2 45.2 80 ;
        RECT 34 75.2 38.8 80 ;
        RECT 27.6 75.2 32.4 80 ;
        RECT 21.2 75.2 26 80 ;
        RECT 14.8 75.2 19.6 80 ;
        RECT 8.4 75.2 13.2 80 ;
        RECT 2 75.2 6.8 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
        RECT 2.65 79.19 5.65 80 ;
    END
    PORT
      LAYER QB ;
        RECT 53.2 0 58 2.4 ;
        RECT 2 24 58 28.8 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER QA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER JA ;
        RECT 53.2 0 58 2.4 ;
        RECT 46.8 0 51.6 2.4 ;
        RECT 40.4 0 45.2 2.4 ;
        RECT 34 0 38.8 2.4 ;
        RECT 27.6 0 32.4 2.4 ;
        RECT 21.2 0 26 2.4 ;
        RECT 14.8 0 19.6 2.4 ;
        RECT 8.4 0 13.2 2.4 ;
        RECT 2 0 6.8 2.4 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END VSUP
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 0 42.6 60 47.4 ;
    END
    PORT
      LAYER QB ;
        RECT 0 17.8 60 22.6 ;
    END
    PORT
      LAYER QB ;
        RECT 0 5.4 60 10.2 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 0 61.2 60 66 ;
    END
    PORT
      LAYER QB ;
        RECT 0 55 60 59.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 0 67.4 60 72.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 48.8 60 53.6 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 0 36.4 60 41.2 ;
    END
    PORT
      LAYER QB ;
        RECT 0 30.2 60 35 ;
    END
    PORT
      LAYER QB ;
        RECT 0 11.6 60 16.4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER JV ;
      RECT 0 0 60 80 ;
    LAYER YS ;
      RECT 0 0 60 80 ;
    LAYER JW ;
      RECT 0 0 60 80 ;
    LAYER QB ;
      RECT 0 0 60 80 ;
    LAYER QA ;
      RECT 0 0 60 80 ;
    LAYER JA ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_IO_SIG_V

MACRO RIIO_EG1D80V_ANACORE_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ANACORE_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 95.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 567.2075 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 54.48 LAYER JA ;
    ANTENNAPARTIALMETALAREA 761.34 LAYER QA ;
    ANTENNAPARTIALMETALAREA 396.54 LAYER QB ;
    ANTENNAPARTIALMETALAREA 188.175 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 12.04192 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 23.04 LAYER JV ;
    ANTENNAPARTIALCUTAREA 54.72 LAYER JW ;
    ANTENNAPARTIALCUTAREA 4.232096 LAYER A2 ;
    ANTENNADIFFAREA 133.0532 LAYER C4 ;
    ANTENNADIFFAREA 133.0532 LAYER C3 ;
    ANTENNADIFFAREA 133.0532 LAYER C5 ;
    ANTENNADIFFAREA 133.0532 LAYER JA ;
    ANTENNADIFFAREA 133.0532 LAYER QA ;
    ANTENNADIFFAREA 133.0532 LAYER QB ;
    ANTENNADIFFAREA 133.0532 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER JA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 24 2 28.8 58 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN VRES3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.735 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 79.654 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 93.78 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.105 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.3648 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 11.75 80 12.25 ;
        RECT 78.15 12.525 80 13.025 ;
        RECT 78.15 13.3 80 13.8 ;
        RECT 78.15 14.075 80 14.575 ;
        RECT 78.15 14.85 80 15.35 ;
      LAYER M2 ;
        RECT 78.15 11.75 80 12.25 ;
        RECT 78.15 12.525 80 13.025 ;
        RECT 78.15 13.3 80 13.8 ;
        RECT 78.15 14.075 80 14.575 ;
        RECT 78.15 14.85 80 15.35 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER JA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER QB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER QA ;
        RECT 77.975 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 78.15 12.05 80 15.05 ;
    END
  END VRES3_B
  PIN VESD0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 24.7745 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 93.505 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 62.855 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 49.35 80 49.85 ;
        RECT 78.15 50.125 80 50.625 ;
        RECT 78.15 50.9 80 51.4 ;
        RECT 78.15 51.675 80 52.175 ;
        RECT 78.15 52.45 80 52.95 ;
      LAYER M2 ;
        RECT 78.15 49.35 80 49.85 ;
        RECT 78.15 50.125 80 50.625 ;
        RECT 78.15 50.9 80 51.4 ;
        RECT 78.15 51.675 80 52.175 ;
        RECT 78.15 52.45 80 52.95 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER JA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER QB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER QA ;
        RECT 77.975 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 78.15 49.65 80 52.65 ;
    END
  END VESD0_B
  PIN VRES0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.235 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 36.0415 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 91.905 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.105 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.099 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.747296 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.6144 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.1664 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 44.65 80 45.15 ;
        RECT 78.15 45.425 80 45.925 ;
        RECT 78.15 46.2 80 46.7 ;
        RECT 78.15 46.975 80 47.475 ;
        RECT 78.15 47.75 80 48.25 ;
      LAYER M2 ;
        RECT 78.15 44.65 80 45.15 ;
        RECT 78.15 45.425 80 45.925 ;
        RECT 78.15 46.2 80 46.7 ;
        RECT 78.15 46.975 80 47.475 ;
        RECT 78.15 47.75 80 48.25 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER JA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER QB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER QA ;
        RECT 77.975 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 78.15 44.95 80 47.95 ;
    END
  END VRES0_B
  PIN VRES1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.235 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 22.887 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 87.235 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 39.95 80 40.45 ;
        RECT 78.15 40.725 80 41.225 ;
        RECT 78.15 41.5 80 42 ;
        RECT 78.15 42.275 80 42.775 ;
        RECT 78.15 43.05 80 43.55 ;
      LAYER M2 ;
        RECT 78.15 39.95 80 40.45 ;
        RECT 78.15 40.725 80 41.225 ;
        RECT 78.15 41.5 80 42 ;
        RECT 78.15 42.275 80 42.775 ;
        RECT 78.15 43.05 80 43.55 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER JA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER QB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER QA ;
        RECT 77.975 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 78.15 40.25 80 43.25 ;
    END
  END VRES1_B
  PIN VESD3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 24.7745 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 93.505 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 62.855 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 7.05 80 7.55 ;
        RECT 78.15 7.825 80 8.325 ;
        RECT 78.15 8.6 80 9.1 ;
        RECT 78.15 9.375 80 9.875 ;
        RECT 78.15 10.15 80 10.65 ;
      LAYER M2 ;
        RECT 78.15 7.05 80 7.55 ;
        RECT 78.15 7.825 80 8.325 ;
        RECT 78.15 8.6 80 9.1 ;
        RECT 78.15 9.375 80 9.875 ;
        RECT 78.15 10.15 80 10.65 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER JA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER QB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER QA ;
        RECT 77.975 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VESD3_B
  PIN VESD2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 21.2495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 96.1675 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.304864 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 21.15 80 21.65 ;
        RECT 78.15 21.925 80 22.425 ;
        RECT 78.15 22.7 80 23.2 ;
        RECT 78.15 23.475 80 23.975 ;
        RECT 78.15 24.25 80 24.75 ;
      LAYER M2 ;
        RECT 78.15 21.15 80 21.65 ;
        RECT 78.15 21.925 80 22.425 ;
        RECT 78.15 22.7 80 23.2 ;
        RECT 78.15 23.475 80 23.975 ;
        RECT 78.15 24.25 80 24.75 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER JA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER QB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER QA ;
        RECT 77.975 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 78.15 21.45 80 24.45 ;
    END
  END VESD2_B
  PIN VRES2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.735 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 21.257 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 85.36 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.747296 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.2624 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 16.45 80 16.95 ;
        RECT 78.15 17.225 80 17.725 ;
        RECT 78.15 18 80 18.5 ;
        RECT 78.15 18.775 80 19.275 ;
        RECT 78.15 19.55 80 20.05 ;
      LAYER M2 ;
        RECT 78.15 16.45 80 16.95 ;
        RECT 78.15 17.225 80 17.725 ;
        RECT 78.15 18 80 18.5 ;
        RECT 78.15 18.775 80 19.275 ;
        RECT 78.15 19.55 80 20.05 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER JA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER QB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER QA ;
        RECT 77.975 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 78.15 16.75 80 19.75 ;
    END
  END VRES2_B
  PIN VESD1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 42.1975 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 98.0425 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.3392 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 35.25 80 35.75 ;
        RECT 78.15 36.025 80 36.525 ;
        RECT 78.15 36.8 80 37.3 ;
        RECT 78.15 37.575 80 38.075 ;
        RECT 78.15 38.35 80 38.85 ;
      LAYER M2 ;
        RECT 78.15 35.25 80 35.75 ;
        RECT 78.15 36.025 80 36.525 ;
        RECT 78.15 36.8 80 37.3 ;
        RECT 78.15 37.575 80 38.075 ;
        RECT 78.15 38.35 80 38.85 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER JA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER QB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER QA ;
        RECT 77.975 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 78.15 35.55 80 38.55 ;
    END
  END VESD1_B
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_ANACORE_H

MACRO RIIO_EG1D80V_ANAIO_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ANAIO_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 95.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 567.2075 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 54.48 LAYER JA ;
    ANTENNAPARTIALMETALAREA 761.34 LAYER QA ;
    ANTENNAPARTIALMETALAREA 396.54 LAYER QB ;
    ANTENNAPARTIALMETALAREA 124.425 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 12.04192 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 23.04 LAYER JV ;
    ANTENNAPARTIALCUTAREA 54.72 LAYER JW ;
    ANTENNAPARTIALCUTAREA 4.905824 LAYER A2 ;
    ANTENNADIFFAREA 148.5876 LAYER C4 ;
    ANTENNADIFFAREA 148.5876 LAYER C3 ;
    ANTENNADIFFAREA 148.5876 LAYER C5 ;
    ANTENNADIFFAREA 148.5876 LAYER JA ;
    ANTENNADIFFAREA 148.5876 LAYER QA ;
    ANTENNADIFFAREA 148.5876 LAYER QB ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER JA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 24 2 28.8 58 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN VRES3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 85.987 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 138.78 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.105 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.099 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.747296 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.6144 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.1664 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 44.65 80 45.15 ;
        RECT 78.15 45.425 80 45.925 ;
        RECT 78.15 46.2 80 46.7 ;
        RECT 78.15 46.975 80 47.475 ;
        RECT 78.15 47.75 80 48.25 ;
      LAYER M2 ;
        RECT 78.15 44.65 80 45.15 ;
        RECT 78.15 45.425 80 45.925 ;
        RECT 78.15 46.2 80 46.7 ;
        RECT 78.15 46.975 80 47.475 ;
        RECT 78.15 47.75 80 48.25 ;
      LAYER C1 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER JA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER QB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER QA ;
        RECT 77.975 44.95 80 47.95 ;
    END
  END VRES3_B
  PIN VESD0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 43.4095 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 138.505 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 62.855 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 7.05 80 7.55 ;
        RECT 78.15 7.825 80 8.325 ;
        RECT 78.15 8.6 80 9.1 ;
        RECT 78.15 9.375 80 9.875 ;
        RECT 78.15 10.15 80 10.65 ;
      LAYER M2 ;
        RECT 78.15 7.05 80 7.55 ;
        RECT 78.15 7.825 80 8.325 ;
        RECT 78.15 8.6 80 9.1 ;
        RECT 78.15 9.375 80 9.875 ;
        RECT 78.15 10.15 80 10.65 ;
      LAYER C1 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER JA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER QB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER QA ;
        RECT 77.975 7.35 80 10.35 ;
    END
  END VESD0_B
  PIN VRES0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.735 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 115.654 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 138.78 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.105 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.3648 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 11.75 80 12.25 ;
        RECT 78.15 12.525 80 13.025 ;
        RECT 78.15 13.3 80 13.8 ;
        RECT 78.15 14.075 80 14.575 ;
        RECT 78.15 14.85 80 15.35 ;
      LAYER M2 ;
        RECT 78.15 11.75 80 12.25 ;
        RECT 78.15 12.525 80 13.025 ;
        RECT 78.15 13.3 80 13.8 ;
        RECT 78.15 14.075 80 14.575 ;
        RECT 78.15 14.85 80 15.35 ;
      LAYER C1 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER JA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER QB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER QA ;
        RECT 77.975 12.05 80 15.05 ;
    END
  END VRES0_B
  PIN VRES1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.86 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 30.257 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 132.235 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.747296 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.2624 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 16.45 80 16.95 ;
        RECT 78.15 17.225 80 17.725 ;
        RECT 78.15 18 80 18.5 ;
        RECT 78.15 18.775 80 19.275 ;
        RECT 78.15 19.55 80 20.05 ;
      LAYER M2 ;
        RECT 78.15 16.45 80 16.95 ;
        RECT 78.15 17.225 80 17.725 ;
        RECT 78.15 18 80 18.5 ;
        RECT 78.15 18.775 80 19.275 ;
        RECT 78.15 19.55 80 20.05 ;
      LAYER C1 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER JA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER QB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER QA ;
        RECT 77.975 16.75 80 19.75 ;
    END
  END VRES1_B
  PIN VESD3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 43.4095 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 138.505 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 62.855 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 3.42792 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 49.35 80 49.85 ;
        RECT 78.15 50.125 80 50.625 ;
        RECT 78.15 50.9 80 51.4 ;
        RECT 78.15 51.675 80 52.175 ;
        RECT 78.15 52.45 80 52.95 ;
      LAYER M2 ;
        RECT 78.15 49.35 80 49.85 ;
        RECT 78.15 50.125 80 50.625 ;
        RECT 78.15 50.9 80 51.4 ;
        RECT 78.15 51.675 80 52.175 ;
        RECT 78.15 52.45 80 52.95 ;
      LAYER C1 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER JA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER QB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER QA ;
        RECT 77.975 49.65 80 52.65 ;
    END
  END VESD3_B
  PIN VESD2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 60.1975 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 143.805 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.3392 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 35.25 80 35.75 ;
        RECT 78.15 36.025 80 36.525 ;
        RECT 78.15 36.8 80 37.3 ;
        RECT 78.15 37.575 80 38.075 ;
        RECT 78.15 38.35 80 38.85 ;
      LAYER M2 ;
        RECT 78.15 35.25 80 35.75 ;
        RECT 78.15 36.025 80 36.525 ;
        RECT 78.15 36.8 80 37.3 ;
        RECT 78.15 37.575 80 38.075 ;
        RECT 78.15 38.35 80 38.85 ;
      LAYER C1 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER JA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER QB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER QA ;
        RECT 77.975 35.55 80 38.55 ;
    END
  END VESD2_B
  PIN VRES2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.235 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 41.522 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 132.235 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 39.95 80 40.45 ;
        RECT 78.15 40.725 80 41.225 ;
        RECT 78.15 41.5 80 42 ;
        RECT 78.15 42.275 80 42.775 ;
        RECT 78.15 43.05 80 43.55 ;
      LAYER M2 ;
        RECT 78.15 39.95 80 40.45 ;
        RECT 78.15 40.725 80 41.225 ;
        RECT 78.15 41.5 80 42 ;
        RECT 78.15 42.275 80 42.775 ;
        RECT 78.15 43.05 80 43.55 ;
      LAYER C1 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER JA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER QB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER QA ;
        RECT 77.975 40.25 80 43.25 ;
    END
  END VRES2_B
  PIN VESD1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 39.8845 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 143.805 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER JA ;
    ANTENNAPARTIALMETALAREA 9.765 LAYER QA ;
    ANTENNAPARTIALMETALAREA 10.29 LAYER QB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 2.913732 LAYER YS ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JV ;
    ANTENNAPARTIALCUTAREA 2.88 LAYER JW ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER JA ;
    ANTENNADIFFAREA 20.425 LAYER QA ;
    ANTENNADIFFAREA 20.425 LAYER QB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 21.15 80 21.65 ;
        RECT 78.15 21.925 80 22.425 ;
        RECT 78.15 22.7 80 23.2 ;
        RECT 78.15 23.475 80 23.975 ;
        RECT 78.15 24.25 80 24.75 ;
      LAYER M2 ;
        RECT 78.15 21.15 80 21.65 ;
        RECT 78.15 21.925 80 22.425 ;
        RECT 78.15 22.7 80 23.2 ;
        RECT 78.15 23.475 80 23.975 ;
        RECT 78.15 24.25 80 24.75 ;
      LAYER C1 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER JA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER QB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER QA ;
        RECT 77.975 21.45 80 24.45 ;
    END
  END VESD1_B
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_ANAIO_H

MACRO RIIO_EG1D80V_BIASPAD_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_BIASPAD_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.25 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 46.875 LAYER C5 ;
    ANTENNAPARTIALCUTAREA 0.894432 LAYER A4 ;
    ANTENNADIFFAREA 3.608 LAYER C4 ;
    ANTENNADIFFAREA 3.608 LAYER C5 ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER C4 ;
        RECT 39.575 0 40.825 60 ;
    END
  END VBIAS
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 567.2075 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER JA ;
    ANTENNAPARTIALMETALAREA 733.44 LAYER QA ;
    ANTENNAPARTIALMETALAREA 391.68 LAYER QB ;
    ANTENNAPARTIALMETALAREA 381.27 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 30.85128 LAYER YS ;
    ANTENNAPARTIALCUTAREA 54.72 LAYER JV ;
    ANTENNAPARTIALCUTAREA 54.72 LAYER JW ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A2 ;
    ANTENNADIFFAREA 148.5876 LAYER C4 ;
    ANTENNADIFFAREA 148.5876 LAYER C3 ;
    ANTENNADIFFAREA 148.5876 LAYER C5 ;
    ANTENNADIFFAREA 148.5876 LAYER JA ;
    ANTENNADIFFAREA 148.5876 LAYER QA ;
    ANTENNADIFFAREA 148.5876 LAYER QB ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_BIASPAD_H

MACRO RIIO_EG1D80V_CUTB2B_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTB2B_H 0 0 ;
  SIZE 80 BY 16 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_l VSS_L!" ;
    PORT
      LAYER QB ;
        RECT 48.8 8.875 53.6 16 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 8.875 72.2 16 ;
    END
  END VSS_L
  PIN VSSIO_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_r VSSIO_R!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 7.125 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 7.125 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 7.125 ;
    END
  END VSSIO_R
  PIN VSS_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_r VSS_R!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 7.125 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 7.125 ;
    END
  END VSS_R
  PIN VSSIO_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_l VSSIO_L!" ;
    PORT
      LAYER QB ;
        RECT 5.4 8.875 10.2 16 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 8.875 22.6 16 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 8.875 47.4 16 ;
    END
  END VSSIO_L
  OBS
    LAYER CA ;
      RECT 0 0 80 16 ;
    LAYER M1 ;
      RECT 0 0 80 16 ;
    LAYER V1 ;
      RECT 0 0 80 16 ;
    LAYER M2 ;
      RECT 0 0 80 16 ;
    LAYER A1 ;
      RECT 0 0 80 16 ;
    LAYER C2 ;
      RECT 0 0 80 16 ;
    LAYER CB ;
      RECT 0 0 80 16 ;
    LAYER JV ;
      RECT 0 0 80 16 ;
    LAYER YS ;
      RECT 0 0 80 16 ;
    LAYER JW ;
      RECT 0 0 80 16 ;
    LAYER QB ;
      RECT 0 0 80 16 ;
    LAYER QA ;
      RECT 0 0 80 16 ;
    LAYER JA ;
      RECT 0 0 80 16 ;
    LAYER AY ;
      RECT 0 0 80 16 ;
    LAYER C1 ;
      RECT 0 0 80 16 ;
    LAYER C5 ;
      RECT 0 0 80 16 ;
    LAYER C4 ;
      RECT 0 0 80 16 ;
    LAYER C3 ;
      RECT 0 0 80 16 ;
    LAYER A4 ;
      RECT 0 0 80 16 ;
    LAYER A3 ;
      RECT 0 0 80 16 ;
    LAYER A2 ;
      RECT 0 0 80 16 ;
  END
END RIIO_EG1D80V_CUTB2B_H

MACRO RIIO_EG1D80V_CUTBIAS_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTBIAS_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 4 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 4 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 4 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 4 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 4 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTBIAS_H

MACRO RIIO_EG1D80V_CUTCOREB2B_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCOREB2B_H 0 0 ;
  SIZE 80 BY 16 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 16 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 16 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 16 ;
    END
  END VSSIO
  PIN VSS_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_r VSS_R!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 7.125 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 7.125 ;
    END
  END VSS_R
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 16 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 16 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 16 ;
    END
  END VDDIO
  PIN VSS_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_l VSS_L!" ;
    PORT
      LAYER QB ;
        RECT 48.8 8.875 53.6 16 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 8.875 72.2 16 ;
    END
  END VSS_L
  OBS
    LAYER CA ;
      RECT 0 0 80 16 ;
    LAYER M1 ;
      RECT 0 0 80 16 ;
    LAYER V1 ;
      RECT 0 0 80 16 ;
    LAYER M2 ;
      RECT 0 0 80 16 ;
    LAYER A1 ;
      RECT 0 0 80 16 ;
    LAYER C2 ;
      RECT 0 0 80 16 ;
    LAYER CB ;
      RECT 0 0 80 16 ;
    LAYER JV ;
      RECT 0 0 80 16 ;
    LAYER YS ;
      RECT 0 0 80 16 ;
    LAYER JW ;
      RECT 0 0 80 16 ;
    LAYER QB ;
      RECT 0 0 80 16 ;
    LAYER QA ;
      RECT 0 0 80 16 ;
    LAYER JA ;
      RECT 0 0 80 16 ;
    LAYER AY ;
      RECT 0 0 80 16 ;
    LAYER C1 ;
      RECT 0 0 80 16 ;
    LAYER C5 ;
      RECT 0 0 80 16 ;
    LAYER C4 ;
      RECT 0 0 80 16 ;
    LAYER C3 ;
      RECT 0 0 80 16 ;
    LAYER A4 ;
      RECT 0 0 80 16 ;
    LAYER A3 ;
      RECT 0 0 80 16 ;
    LAYER A2 ;
      RECT 0 0 80 16 ;
  END
END RIIO_EG1D80V_CUTCOREB2B_H

MACRO RIIO_EG1D80V_CUTCOREPWR_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCOREPWR_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 4 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 4 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 4 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 4 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTCOREPWR_H

MACRO RIIO_EG1D80V_CUTCORE_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCORE_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 4 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 4 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 4 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTCORE_H

MACRO RIIO_EG1D80V_CUTIOB2B_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIOB2B_H 0 0 ;
  SIZE 80 BY 16 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_l VSSIO_L!" ;
    PORT
      LAYER QB ;
        RECT 5.4 8.875 10.2 16 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 8.875 22.6 16 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 8.875 47.4 16 ;
    END
  END VSSIO_L
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 16 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 16 ;
    END
  END VDD
  PIN VSSIO_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_r VSSIO_R!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 7.125 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 7.125 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 7.125 ;
    END
  END VSSIO_R
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 16 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 16 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 16 ;
    LAYER M1 ;
      RECT 0 0 80 16 ;
    LAYER V1 ;
      RECT 0 0 80 16 ;
    LAYER M2 ;
      RECT 0 0 80 16 ;
    LAYER A1 ;
      RECT 0 0 80 16 ;
    LAYER C2 ;
      RECT 0 0 80 16 ;
    LAYER CB ;
      RECT 0 0 80 16 ;
    LAYER JV ;
      RECT 0 0 80 16 ;
    LAYER YS ;
      RECT 0 0 80 16 ;
    LAYER JW ;
      RECT 0 0 80 16 ;
    LAYER QB ;
      RECT 0 0 80 16 ;
    LAYER QA ;
      RECT 0 0 80 16 ;
    LAYER JA ;
      RECT 0 0 80 16 ;
    LAYER AY ;
      RECT 0 0 80 16 ;
    LAYER C1 ;
      RECT 0 0 80 16 ;
    LAYER C5 ;
      RECT 0 0 80 16 ;
    LAYER C4 ;
      RECT 0 0 80 16 ;
    LAYER C3 ;
      RECT 0 0 80 16 ;
    LAYER A4 ;
      RECT 0 0 80 16 ;
    LAYER A3 ;
      RECT 0 0 80 16 ;
    LAYER A2 ;
      RECT 0 0 80 16 ;
  END
END RIIO_EG1D80V_CUTIOB2B_H

MACRO RIIO_EG1D80V_CUTIOPWR_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIOPWR_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 4 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 4 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 4 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTIOPWR_H

MACRO RIIO_EG1D80V_CUTIO_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIO_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 4 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 4 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTIO_H

MACRO RIIO_EG1D80V_CUTPWR_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTPWR_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 4 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 4 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTPWR_H

MACRO RIIO_EG1D80V_CUT_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUT_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUT_H

MACRO RIIO_EG1D80V_FILL16B2B_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL16B2B_H 0 0 ;
  SIZE 80 BY 16 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 16 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 16 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 16 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 16 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 16 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 16 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 16 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 16 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 16 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 16 ;
    LAYER M1 ;
      RECT 0 0 80 16 ;
    LAYER V1 ;
      RECT 0 0 80 16 ;
    LAYER M2 ;
      RECT 0 0 80 16 ;
    LAYER A1 ;
      RECT 0 0 80 16 ;
    LAYER C2 ;
      RECT 0 0 80 16 ;
    LAYER CB ;
      RECT 0 0 80 16 ;
    LAYER JV ;
      RECT 0 0 80 16 ;
    LAYER YS ;
      RECT 0 0 80 16 ;
    LAYER JW ;
      RECT 0 0 80 16 ;
    LAYER QB ;
      RECT 0 0 80 16 ;
    LAYER QA ;
      RECT 0 0 80 16 ;
    LAYER JA ;
      RECT 0 0 80 16 ;
    LAYER AY ;
      RECT 0 0 80 16 ;
    LAYER C1 ;
      RECT 0 0 80 16 ;
    LAYER C5 ;
      RECT 0 0 80 16 ;
    LAYER C4 ;
      RECT 0 0 80 16 ;
    LAYER C3 ;
      RECT 0 0 80 16 ;
    LAYER A4 ;
      RECT 0 0 80 16 ;
    LAYER A3 ;
      RECT 0 0 80 16 ;
    LAYER A2 ;
      RECT 0 0 80 16 ;
  END
END RIIO_EG1D80V_FILL16B2B_H

MACRO RIIO_EG1D80V_FILL16_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL16_H 0 0 ;
  SIZE 80 BY 16 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 16 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 16 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 16 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 16 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 16 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 16 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 16 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 16 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 16 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 16 ;
    LAYER M1 ;
      RECT 0 0 80 16 ;
    LAYER V1 ;
      RECT 0 0 80 16 ;
    LAYER M2 ;
      RECT 0 0 80 16 ;
    LAYER A1 ;
      RECT 0 0 80 16 ;
    LAYER C2 ;
      RECT 0 0 80 16 ;
    LAYER CB ;
      RECT 0 0 80 16 ;
    LAYER JV ;
      RECT 0 0 80 16 ;
    LAYER YS ;
      RECT 0 0 80 16 ;
    LAYER JW ;
      RECT 0 0 80 16 ;
    LAYER QB ;
      RECT 0 0 80 16 ;
    LAYER QA ;
      RECT 0 0 80 16 ;
    LAYER JA ;
      RECT 0 0 80 16 ;
    LAYER AY ;
      RECT 0 0 80 16 ;
    LAYER C1 ;
      RECT 0 0 80 16 ;
    LAYER C5 ;
      RECT 0 0 80 16 ;
    LAYER C4 ;
      RECT 0 0 80 16 ;
    LAYER C3 ;
      RECT 0 0 80 16 ;
    LAYER A4 ;
      RECT 0 0 80 16 ;
    LAYER A3 ;
      RECT 0 0 80 16 ;
    LAYER A2 ;
      RECT 0 0 80 16 ;
  END
END RIIO_EG1D80V_FILL16_H

MACRO RIIO_EG1D80V_FILL1_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL1_H 0 0 ;
  SIZE 80 BY 1 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 1 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 1 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 1 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 1 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 1 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 1 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 1 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 1 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 1 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 1 ;
    LAYER M1 ;
      RECT 0 0 80 1 ;
    LAYER V1 ;
      RECT 0 0 80 1 ;
    LAYER M2 ;
      RECT 0 0 80 1 ;
    LAYER A1 ;
      RECT 0 0 80 1 ;
    LAYER C2 ;
      RECT 0 0 80 1 ;
    LAYER CB ;
      RECT 0 0 80 1 ;
    LAYER JV ;
      RECT 0 0 80 1 ;
    LAYER YS ;
      RECT 0 0 80 1 ;
    LAYER JW ;
      RECT 0 0 80 1 ;
    LAYER QB ;
      RECT 0 0 80 1 ;
    LAYER QA ;
      RECT 0 0 80 1 ;
    LAYER JA ;
      RECT 0 0 80 1 ;
    LAYER AY ;
      RECT 0 0 80 1 ;
    LAYER C1 ;
      RECT 0 0 80 1 ;
    LAYER C5 ;
      RECT 0 0 80 1 ;
    LAYER C4 ;
      RECT 0 0 80 1 ;
    LAYER C3 ;
      RECT 0 0 80 1 ;
    LAYER A4 ;
      RECT 0 0 80 1 ;
    LAYER A3 ;
      RECT 0 0 80 1 ;
    LAYER A2 ;
      RECT 0 0 80 1 ;
  END
END RIIO_EG1D80V_FILL1_H

MACRO RIIO_EG1D80V_FILL2_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL2_H 0 0 ;
  SIZE 80 BY 2 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 2 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 2 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 2 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 2 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 2 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 2 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 2 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 2 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 80 2 ;
    LAYER M1 ;
      RECT 0 0 80 2 ;
    LAYER V1 ;
      RECT 0 0 80 2 ;
    LAYER M2 ;
      RECT 0 0 80 2 ;
    LAYER A1 ;
      RECT 0 0 80 2 ;
    LAYER C2 ;
      RECT 0 0 80 2 ;
    LAYER CB ;
      RECT 0 0 80 2 ;
    LAYER JV ;
      RECT 0 0 80 2 ;
    LAYER YS ;
      RECT 0 0 80 2 ;
    LAYER JW ;
      RECT 0 0 80 2 ;
    LAYER QB ;
      RECT 0 0 80 2 ;
    LAYER QA ;
      RECT 0 0 80 2 ;
    LAYER JA ;
      RECT 0 0 80 2 ;
    LAYER AY ;
      RECT 0 0 80 2 ;
    LAYER C1 ;
      RECT 0 0 80 2 ;
    LAYER C5 ;
      RECT 0 0 80 2 ;
    LAYER C4 ;
      RECT 0 0 80 2 ;
    LAYER C3 ;
      RECT 0 0 80 2 ;
    LAYER A4 ;
      RECT 0 0 80 2 ;
    LAYER A3 ;
      RECT 0 0 80 2 ;
    LAYER A2 ;
      RECT 0 0 80 2 ;
  END
END RIIO_EG1D80V_FILL2_H

MACRO RIIO_EG1D80V_FILL32_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL32_H 0 0 ;
  SIZE 80 BY 32 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 32 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 32 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 32 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 32 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 32 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 32 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 32 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 32 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 32 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 32 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 32 ;
    LAYER M1 ;
      RECT 0 0 80 32 ;
    LAYER V1 ;
      RECT 0 0 80 32 ;
    LAYER M2 ;
      RECT 0 0 80 32 ;
    LAYER A1 ;
      RECT 0 0 80 32 ;
    LAYER C2 ;
      RECT 0 0 80 32 ;
    LAYER CB ;
      RECT 0 0 80 32 ;
    LAYER JV ;
      RECT 0 0 80 32 ;
    LAYER YS ;
      RECT 0 0 80 32 ;
    LAYER JW ;
      RECT 0 0 80 32 ;
    LAYER QB ;
      RECT 0 0 80 32 ;
    LAYER QA ;
      RECT 0 0 80 32 ;
    LAYER JA ;
      RECT 0 0 80 32 ;
    LAYER AY ;
      RECT 0 0 80 32 ;
    LAYER C1 ;
      RECT 0 0 80 32 ;
    LAYER C5 ;
      RECT 0 0 80 32 ;
    LAYER C4 ;
      RECT 0 0 80 32 ;
    LAYER C3 ;
      RECT 0 0 80 32 ;
    LAYER A4 ;
      RECT 0 0 80 32 ;
    LAYER A3 ;
      RECT 0 0 80 32 ;
    LAYER A2 ;
      RECT 0 0 80 32 ;
  END
END RIIO_EG1D80V_FILL32_H

MACRO RIIO_EG1D80V_FILL4_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL4_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 4 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 4 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 4 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 4 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 4 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 4 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_FILL4_H

MACRO RIIO_EG1D80V_FILL8_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL8_H 0 0 ;
  SIZE 80 BY 8 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 8 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 8 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 8 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 8 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 8 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 8 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 8 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 8 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 8 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 8 ;
    LAYER M1 ;
      RECT 0 0 80 8 ;
    LAYER V1 ;
      RECT 0 0 80 8 ;
    LAYER M2 ;
      RECT 0 0 80 8 ;
    LAYER A1 ;
      RECT 0 0 80 8 ;
    LAYER C2 ;
      RECT 0 0 80 8 ;
    LAYER CB ;
      RECT 0 0 80 8 ;
    LAYER JV ;
      RECT 0 0 80 8 ;
    LAYER YS ;
      RECT 0 0 80 8 ;
    LAYER JW ;
      RECT 0 0 80 8 ;
    LAYER QB ;
      RECT 0 0 80 8 ;
    LAYER QA ;
      RECT 0 0 80 8 ;
    LAYER JA ;
      RECT 0 0 80 8 ;
    LAYER AY ;
      RECT 0 0 80 8 ;
    LAYER C1 ;
      RECT 0 0 80 8 ;
    LAYER C5 ;
      RECT 0 0 80 8 ;
    LAYER C4 ;
      RECT 0 0 80 8 ;
    LAYER C3 ;
      RECT 0 0 80 8 ;
    LAYER A4 ;
      RECT 0 0 80 8 ;
    LAYER A3 ;
      RECT 0 0 80 8 ;
    LAYER A2 ;
      RECT 0 0 80 8 ;
  END
END RIIO_EG1D80V_FILL8_H

MACRO RIIO_EG1D80V_POR_IO_V1D0_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_POR_IO_V1D0_H 0 0 ;
  SIZE 80 BY 8 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER C3 ;
        RECT 37.075 0 39.575 8 ;
    END
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 8 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 8 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 8 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER C3 ;
        RECT 70.825 0 73.325 8 ;
    END
    PORT
      LAYER QB ;
        RECT 55 0 59.8 8 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER C3 ;
        RECT 74.575 0 77.075 8 ;
    END
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 8 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 8 ;
    END
  END VSS
  PIN VDDIO_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio_por VDDIO_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 33.325 2.625 80 3.125 ;
    END
  END VDDIO_POR
  PIN POR_N_CORE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3375 LAYER C2 ;
    ANTENNADIFFAREA 0.2453 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.5 5.625 80 6.125 ;
    END
  END POR_N_CORE_O
  PIN VDD_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd_por VDD_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 70.825 4.125 80 4.625 ;
    END
  END VDD_POR
  PIN VSSIO_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_por VSSIO_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 33.325 1.875 80 2.375 ;
    END
  END VSSIO_POR
  PIN VSS_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_por VSS_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 70.825 4.875 80 5.375 ;
    END
  END VSS_POR
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 8 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 8 ;
      LAYER C3 ;
        RECT 33.325 0 35.825 8 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 8 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 8 ;
    LAYER M1 ;
      RECT 0 0 80 8 ;
    LAYER V1 ;
      RECT 0 0 80 8 ;
    LAYER M2 ;
      RECT 0 0 80 8 ;
    LAYER A1 ;
      RECT 0 0 80 8 ;
    LAYER C2 ;
      RECT 0 0 80 8 ;
    LAYER CB ;
      RECT 0 0 80 8 ;
    LAYER JV ;
      RECT 0 0 80 8 ;
    LAYER YS ;
      RECT 0 0 80 8 ;
    LAYER JW ;
      RECT 0 0 80 8 ;
    LAYER QB ;
      RECT 0 0 80 8 ;
    LAYER QA ;
      RECT 0 0 80 8 ;
    LAYER JA ;
      RECT 0 0 80 8 ;
    LAYER AY ;
      RECT 0 0 80 8 ;
    LAYER C1 ;
      RECT 0 0 80 8 ;
    LAYER C5 ;
      RECT 0 0 80 8 ;
    LAYER C4 ;
      RECT 0 0 80 8 ;
    LAYER C3 ;
      RECT 0 0 80 8 ;
    LAYER A4 ;
      RECT 0 0 80 8 ;
    LAYER A3 ;
      RECT 0 0 80 8 ;
    LAYER A2 ;
      RECT 0 0 80 8 ;
  END
END RIIO_EG1D80V_POR_IO_V1D0_H

MACRO RIIO_EG1D80V_RAILSHORT_GND_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_GND_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 4 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 4 ;
    END
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 4 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 4 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 4 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_RAILSHORT_GND_H

MACRO RIIO_EG1D80V_RAILSHORT_PG_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_PG_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 4 ;
    END
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 4 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 4 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 55 0 59.8 4 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 4 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_RAILSHORT_PG_H

MACRO RIIO_EG1D80V_RAILSHORT_PWR_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_PWR_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 4 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 4 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 4 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 4 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 4 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 4 ;
    END
    PORT
      LAYER QB ;
        RECT 55 0 59.8 4 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 4 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER JV ;
      RECT 0 0 80 4 ;
    LAYER YS ;
      RECT 0 0 80 4 ;
    LAYER JW ;
      RECT 0 0 80 4 ;
    LAYER QB ;
      RECT 0 0 80 4 ;
    LAYER QA ;
      RECT 0 0 80 4 ;
    LAYER JA ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_RAILSHORT_PWR_H

MACRO RIIO_EG1D80V_VDD04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDD04_H

MACRO RIIO_EG1D80V_VDDIOX_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDIOX_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDDIOX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddiox VDDIOX!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
    END
  END VDDIOX
  PIN VSSIOX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssiox VSSIOX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSSIOX
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDIOX_H

MACRO RIIO_EG1D80V_VDDIO_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDIO_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDIO_H

MACRO RIIO_EG1D80V_VDDQ04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VDDQ
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDQ04_H

MACRO RIIO_EG1D80V_VDDQ_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VDDQ
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDQ_HVT_H

MACRO RIIO_EG1D80V_VDDQ_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VDDQ
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDQ_RVT_H

MACRO RIIO_EG1D80V_VDDX04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
        RECT 78.15 51.25 80 53.75 ;
        RECT 78.15 55 80 57.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
        RECT 78.15 51.25 80 53.75 ;
        RECT 78.15 55 80 57.5 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
        RECT 79.19 51.088 80 51.588 ;
        RECT 79.19 51.863 80 52.363 ;
        RECT 79.19 52.638 80 53.138 ;
        RECT 79.19 53.413 80 53.913 ;
        RECT 79.19 54.838 80 55.338 ;
        RECT 79.19 55.613 80 56.113 ;
        RECT 79.19 56.388 80 56.888 ;
        RECT 79.19 57.163 80 57.663 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
        RECT 79.19 47.338 80 50.163 ;
        RECT 79.19 51.088 80 53.913 ;
        RECT 79.19 54.838 80 57.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
        RECT 79.19 51.088 80 51.588 ;
        RECT 79.19 51.863 80 52.363 ;
        RECT 79.19 52.638 80 53.138 ;
        RECT 79.19 53.413 80 53.913 ;
        RECT 79.19 54.838 80 55.338 ;
        RECT 79.19 55.613 80 56.113 ;
        RECT 79.19 56.388 80 56.888 ;
        RECT 79.19 57.163 80 57.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 2.5 80 5 ;
        RECT 78.15 6.25 80 8.75 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 2.5 80 5 ;
        RECT 78.15 6.25 80 8.75 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER M2 ;
        RECT 79.19 2.338 80 2.838 ;
        RECT 79.19 3.113 80 3.613 ;
        RECT 79.19 3.888 80 4.388 ;
        RECT 79.19 4.663 80 5.163 ;
        RECT 79.19 6.088 80 6.588 ;
        RECT 79.19 6.863 80 7.363 ;
        RECT 79.19 7.638 80 8.138 ;
        RECT 79.19 8.413 80 8.913 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER C1 ;
        RECT 79.19 2.338 80 5.163 ;
        RECT 79.19 6.088 80 8.913 ;
        RECT 79.19 9.838 80 12.663 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 2.338 80 2.838 ;
        RECT 79.19 3.113 80 3.613 ;
        RECT 79.19 3.888 80 4.388 ;
        RECT 79.19 4.663 80 5.163 ;
        RECT 79.19 6.088 80 6.588 ;
        RECT 79.19 6.863 80 7.363 ;
        RECT 79.19 7.638 80 8.138 ;
        RECT 79.19 8.413 80 8.913 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
    END
  END VSSX
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDX04_H

MACRO RIIO_EG1D80V_VDDX_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDX_HVT_H

MACRO RIIO_EG1D80V_VDDX_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDX_RVT_H

MACRO RIIO_EG1D80V_VDD_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDD_HVT_H

MACRO RIIO_EG1D80V_VDD_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDD_RVT_H

MACRO RIIO_EG1D80V_VNWINT_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNWINT_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VNWINT_HVT_H

MACRO RIIO_EG1D80V_VNWINT_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNWINT_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VNWINT_RVT_H

MACRO RIIO_EG1D80V_VNW_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNW_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VNW_H

MACRO RIIO_EG1D80V_VPWINT_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPWINT_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VPWINT_HVT_H

MACRO RIIO_EG1D80V_VPWINT_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPWINT_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VPWINT_RVT_H

MACRO RIIO_EG1D80V_VPW_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPW_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VPW_H

MACRO RIIO_EG1D80V_VSS04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSS04_H

MACRO RIIO_EG1D80V_VSSIOX_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSIOX_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VSSIOX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssiox VSSIOX!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.153 40.25 80.003 43.25 ;
        RECT 78.153 44.95 80.003 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.153 40.25 80.003 43.25 ;
        RECT 78.153 44.95 80.003 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
        RECT 78.15 51.251 80 53.751 ;
        RECT 78.15 55.001 80 57.501 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
        RECT 78.15 51.251 80 53.751 ;
        RECT 78.15 55.001 80 57.501 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
        RECT 79.19 47.338 80 50.163 ;
        RECT 79.19 51.089 80 53.914 ;
        RECT 79.19 54.839 80 57.664 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
        RECT 79.19 51.089 80 51.589 ;
        RECT 79.19 51.864 80 52.364 ;
        RECT 79.19 52.639 80 53.139 ;
        RECT 79.19 53.414 80 53.914 ;
        RECT 79.19 54.839 80 55.339 ;
        RECT 79.19 55.614 80 56.114 ;
        RECT 79.19 56.389 80 56.889 ;
        RECT 79.19 57.164 80 57.664 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
        RECT 79.19 51.089 80 51.589 ;
        RECT 79.19 51.864 80 52.364 ;
        RECT 79.19 52.639 80 53.139 ;
        RECT 79.19 53.414 80 53.914 ;
        RECT 79.19 54.839 80 55.339 ;
        RECT 79.19 55.614 80 56.114 ;
        RECT 79.19 56.389 80 56.889 ;
        RECT 79.19 57.164 80 57.664 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.153 12.05 80.003 15.05 ;
        RECT 78.153 16.75 80.003 19.75 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.153 12.05 80.003 15.05 ;
        RECT 78.153 16.75 80.003 19.75 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 2.499 80 4.999 ;
        RECT 78.15 6.25 80 8.75 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 2.499 80 4.999 ;
        RECT 78.15 6.25 80 8.75 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 2.337 80 5.162 ;
        RECT 79.19 6.088 80 8.913 ;
        RECT 79.19 9.838 80 12.663 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 2.337 80 2.837 ;
        RECT 79.19 3.112 80 3.612 ;
        RECT 79.19 3.887 80 4.387 ;
        RECT 79.19 4.662 80 5.162 ;
        RECT 79.19 6.088 80 6.588 ;
        RECT 79.19 6.863 80 7.363 ;
        RECT 79.19 7.638 80 8.138 ;
        RECT 79.19 8.413 80 8.913 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 2.337 80 2.837 ;
        RECT 79.19 3.112 80 3.612 ;
        RECT 79.19 3.887 80 4.387 ;
        RECT 79.19 4.662 80 5.162 ;
        RECT 79.19 6.088 80 6.588 ;
        RECT 79.19 6.863 80 7.363 ;
        RECT 79.19 7.638 80 8.138 ;
        RECT 79.19 8.413 80 8.913 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
  END VSSIOX
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDDIOX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddiox VDDIOX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
    END
  END VDDIOX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSIOX_H

MACRO RIIO_EG1D80V_VSSIO_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSIO_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSIO_H

MACRO RIIO_EG1D80V_VSSQ04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSQ04_H

MACRO RIIO_EG1D80V_VSSQ_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDQ
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSQ_HVT_H

MACRO RIIO_EG1D80V_VSSQ_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDQ
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSQ_RVT_H

MACRO RIIO_EG1D80V_VSSX04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
        RECT 78.15 51.25 80 53.75 ;
        RECT 78.15 55 80 57.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
        RECT 78.15 51.25 80 53.75 ;
        RECT 78.15 55 80 57.5 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
        RECT 79.19 51.088 80 51.588 ;
        RECT 79.19 51.863 80 52.363 ;
        RECT 79.19 52.638 80 53.138 ;
        RECT 79.19 53.413 80 53.913 ;
        RECT 79.19 54.838 80 55.338 ;
        RECT 79.19 55.613 80 56.113 ;
        RECT 79.19 56.388 80 56.888 ;
        RECT 79.19 57.163 80 57.663 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
        RECT 79.19 51.088 80 51.588 ;
        RECT 79.19 51.863 80 52.363 ;
        RECT 79.19 52.638 80 53.138 ;
        RECT 79.19 53.413 80 53.913 ;
        RECT 79.19 54.838 80 55.338 ;
        RECT 79.19 55.613 80 56.113 ;
        RECT 79.19 56.388 80 56.888 ;
        RECT 79.19 57.163 80 57.663 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
        RECT 79.19 47.338 80 50.163 ;
        RECT 79.19 51.088 80 53.913 ;
        RECT 79.19 54.838 80 57.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 2.5 80 5 ;
        RECT 78.15 6.25 80 8.75 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 2.5 80 5 ;
        RECT 78.15 6.25 80 8.75 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER M1 ;
        RECT 79.19 2.338 80 2.838 ;
        RECT 79.19 3.113 80 3.613 ;
        RECT 79.19 3.888 80 4.388 ;
        RECT 79.19 4.663 80 5.163 ;
        RECT 79.19 6.088 80 6.588 ;
        RECT 79.19 6.863 80 7.363 ;
        RECT 79.19 7.638 80 8.138 ;
        RECT 79.19 8.413 80 8.913 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 2.338 80 2.838 ;
        RECT 79.19 3.113 80 3.613 ;
        RECT 79.19 3.888 80 4.388 ;
        RECT 79.19 4.663 80 5.163 ;
        RECT 79.19 6.088 80 6.588 ;
        RECT 79.19 6.863 80 7.363 ;
        RECT 79.19 7.638 80 8.138 ;
        RECT 79.19 8.413 80 8.913 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER C1 ;
        RECT 79.19 2.338 80 5.163 ;
        RECT 79.19 6.088 80 8.913 ;
        RECT 79.19 9.838 80 12.663 ;
        RECT 79.19 17.338 80 20.163 ;
    END
  END VSSX
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSX04_H

MACRO RIIO_EG1D80V_VSSX_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
        RECT 78.15 51.25 80 53.75 ;
        RECT 78.15 55 80 57.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
        RECT 78.15 51.25 80 53.75 ;
        RECT 78.15 55 80 57.5 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
        RECT 79.19 47.338 80 50.163 ;
        RECT 79.19 51.088 80 53.913 ;
        RECT 79.19 54.838 80 57.663 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
        RECT 79.19 51.088 80 51.588 ;
        RECT 79.19 51.863 80 52.363 ;
        RECT 79.19 52.638 80 53.138 ;
        RECT 79.19 53.413 80 53.913 ;
        RECT 79.19 54.838 80 55.338 ;
        RECT 79.19 55.613 80 56.113 ;
        RECT 79.19 56.388 80 56.888 ;
        RECT 79.19 57.163 80 57.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
        RECT 79.19 51.088 80 51.588 ;
        RECT 79.19 51.863 80 52.363 ;
        RECT 79.19 52.638 80 53.138 ;
        RECT 79.19 53.413 80 53.913 ;
        RECT 79.19 54.838 80 55.338 ;
        RECT 79.19 55.613 80 56.113 ;
        RECT 79.19 56.388 80 56.888 ;
        RECT 79.19 57.163 80 57.663 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 2.5 80 5 ;
        RECT 78.15 6.25 80 8.75 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 2.5 80 5 ;
        RECT 78.15 6.25 80 8.75 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 2.338 80 5.163 ;
        RECT 79.19 6.088 80 8.913 ;
        RECT 79.19 9.838 80 12.663 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 2.338 80 2.838 ;
        RECT 79.19 3.113 80 3.613 ;
        RECT 79.19 3.888 80 4.388 ;
        RECT 79.19 4.663 80 5.163 ;
        RECT 79.19 6.088 80 6.588 ;
        RECT 79.19 6.863 80 7.363 ;
        RECT 79.19 7.638 80 8.138 ;
        RECT 79.19 8.413 80 8.913 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 2.338 80 2.838 ;
        RECT 79.19 3.113 80 3.613 ;
        RECT 79.19 3.888 80 4.388 ;
        RECT 79.19 4.663 80 5.163 ;
        RECT 79.19 6.088 80 6.588 ;
        RECT 79.19 6.863 80 7.363 ;
        RECT 79.19 7.638 80 8.138 ;
        RECT 79.19 8.413 80 8.913 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSX_HVT_H

MACRO RIIO_EG1D80V_VSSX_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
        RECT 78.15 51.25 80 53.75 ;
        RECT 78.15 55 80 57.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
        RECT 78.15 47.5 80 50 ;
        RECT 78.15 51.25 80 53.75 ;
        RECT 78.15 55 80 57.5 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
        RECT 79.19 47.338 80 50.163 ;
        RECT 79.19 51.088 80 53.913 ;
        RECT 79.19 54.838 80 57.663 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
        RECT 79.19 51.088 80 51.588 ;
        RECT 79.19 51.863 80 52.363 ;
        RECT 79.19 52.638 80 53.138 ;
        RECT 79.19 53.413 80 53.913 ;
        RECT 79.19 54.838 80 55.338 ;
        RECT 79.19 55.613 80 56.113 ;
        RECT 79.19 56.388 80 56.888 ;
        RECT 79.19 57.163 80 57.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
        RECT 79.19 51.088 80 51.588 ;
        RECT 79.19 51.863 80 52.363 ;
        RECT 79.19 52.638 80 53.138 ;
        RECT 79.19 53.413 80 53.913 ;
        RECT 79.19 54.838 80 55.338 ;
        RECT 79.19 55.613 80 56.113 ;
        RECT 79.19 56.388 80 56.888 ;
        RECT 79.19 57.163 80 57.663 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.075 80 15.075 ;
        RECT 78.15 16.775 80 19.775 ;
      LAYER C3 ;
        RECT 78.15 2.5 80 5 ;
        RECT 78.15 6.25 80 8.75 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 2.5 80 5 ;
        RECT 78.15 6.25 80 8.75 ;
        RECT 78.15 10 80 12.5 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 2.338 80 5.163 ;
        RECT 79.19 6.088 80 8.913 ;
        RECT 79.19 9.838 80 12.663 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 2.338 80 2.838 ;
        RECT 79.19 3.113 80 3.613 ;
        RECT 79.19 3.888 80 4.388 ;
        RECT 79.19 4.663 80 5.163 ;
        RECT 79.19 6.088 80 6.588 ;
        RECT 79.19 6.863 80 7.363 ;
        RECT 79.19 7.638 80 8.138 ;
        RECT 79.19 8.413 80 8.913 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 2.338 80 2.838 ;
        RECT 79.19 3.113 80 3.613 ;
        RECT 79.19 3.888 80 4.388 ;
        RECT 79.19 4.663 80 5.163 ;
        RECT 79.19 6.088 80 6.588 ;
        RECT 79.19 6.863 80 7.363 ;
        RECT 79.19 7.638 80 8.138 ;
        RECT 79.19 8.413 80 8.913 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER QB ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER JA ;
        RECT 75.2 27.6 80 32.4 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER QB ;
        RECT 75.2 27.6 80 32.4 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSX_RVT_H

MACRO RIIO_EG1D80V_VSS_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSS_HVT_H

MACRO RIIO_EG1D80V_VSS_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
    PORT
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
    END
    PORT
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
    END
    PORT
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
    END
    PORT
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
    END
    PORT
      CLASS CORE ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSS_RVT_H

MACRO RIIO_EG1D80V_VSUP_CORE_GND_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_GND_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VSUP
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_CORE_GND_H

MACRO RIIO_EG1D80V_VSUP_CORE_PWR_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_PWR_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VSUP
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_CORE_PWR_H

MACRO RIIO_EG1D80V_VSUP_CORE_SIG_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_SIG_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.633 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1122.47 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 610.45 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 610.4525 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1151.7 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 660.48 LAYER JA ;
    ANTENNAPARTIALMETALAREA 357.12 LAYER QA ;
    ANTENNAPARTIALMETALAREA 660.48 LAYER QB ;
    ANTENNAPARTIALMETALAREA 4.554 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 2.392896 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 1.792 LAYER AY ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 46.27692 LAYER YS ;
    ANTENNAPARTIALCUTAREA 106.56 LAYER JV ;
    ANTENNAPARTIALCUTAREA 106.56 LAYER JW ;
    ANTENNAPARTIALCUTAREA 1.92 LAYER V1 ;
    ANTENNADIFFAREA 133.0532 LAYER C4 ;
    ANTENNADIFFAREA 133.0532 LAYER C3 ;
    ANTENNADIFFAREA 133.0532 LAYER C5 ;
    ANTENNADIFFAREA 133.0532 LAYER JA ;
    ANTENNADIFFAREA 133.0532 LAYER QA ;
    ANTENNADIFFAREA 133.0532 LAYER QB ;
    ANTENNADIFFAREA 133.0532 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
        RECT 79.19 54.35 80 57.35 ;
    END
  END VSUP
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_CORE_SIG_H

MACRO RIIO_EG1D80V_VSUP_IO_GND_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_GND_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VSUP
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_IO_GND_H

MACRO RIIO_EG1D80V_VSUP_IO_PWR_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_PWR_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER QB ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER QB ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER QA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER JA ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER QB ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER QA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER JA ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER QB ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER QA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER JA ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER QB ;
        RECT 0 2 2.4 6.8 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER QA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER JA ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER QA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER JA ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER QA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER JA ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VSUP
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_IO_PWR_H

MACRO RIIO_EG1D80V_VSUP_IO_SIG_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_SIG_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.633 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1151.7 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 747.95 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 611.5625 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1151.7 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 648.96 LAYER JA ;
    ANTENNAPARTIALMETALAREA 364.8 LAYER QA ;
    ANTENNAPARTIALMETALAREA 660.48 LAYER QB ;
    ANTENNAPARTIALMETALAREA 4.554 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 2.392896 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 1.792 LAYER AY ;
    ANTENNAPARTIALCUTAREA 26.515456 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 46.27692 LAYER YS ;
    ANTENNAPARTIALCUTAREA 106.56 LAYER JV ;
    ANTENNAPARTIALCUTAREA 106.56 LAYER JW ;
    ANTENNAPARTIALCUTAREA 1.92 LAYER V1 ;
    ANTENNADIFFAREA 148.5876 LAYER C4 ;
    ANTENNADIFFAREA 148.5876 LAYER C3 ;
    ANTENNADIFFAREA 148.5876 LAYER C5 ;
    ANTENNADIFFAREA 148.5876 LAYER JA ;
    ANTENNADIFFAREA 148.5876 LAYER QA ;
    ANTENNADIFFAREA 148.5876 LAYER QB ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER QB ;
        RECT 24 2 28.8 58 ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER QA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER JA ;
        RECT 0 2 2.4 6.8 ;
        RECT 0 8.4 2.4 13.2 ;
        RECT 0 14.8 2.4 19.6 ;
        RECT 0 21.2 2.4 26 ;
        RECT 0 27.6 2.4 32.4 ;
        RECT 0 34 2.4 38.8 ;
        RECT 0 40.4 2.4 45.2 ;
        RECT 0 46.8 2.4 51.6 ;
        RECT 0 53.2 2.4 58 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER QB ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER QA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER JA ;
        RECT 75.2 2 80 6.8 ;
        RECT 75.2 8.4 80 13.2 ;
        RECT 75.2 14.8 80 19.6 ;
        RECT 75.2 21.2 80 26 ;
        RECT 75.2 27.6 80 32.4 ;
        RECT 75.2 34 80 38.8 ;
        RECT 75.2 40.4 80 45.2 ;
        RECT 75.2 46.8 80 51.6 ;
        RECT 75.2 53.2 80 58 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
        RECT 79.19 54.35 80 57.35 ;
    END
  END VSUP
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER QB ;
        RECT 48.8 0 53.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 67.4 0 72.2 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER QB ;
        RECT 11.6 0 16.4 60 ;
    END
    PORT
      LAYER QB ;
        RECT 30.2 0 35 60 ;
    END
    PORT
      LAYER QB ;
        RECT 36.4 0 41.2 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER QB ;
        RECT 5.4 0 10.2 60 ;
    END
    PORT
      LAYER QB ;
        RECT 17.8 0 22.6 60 ;
    END
    PORT
      LAYER QB ;
        RECT 42.6 0 47.4 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER QB ;
        RECT 55 0 59.8 60 ;
    END
    PORT
      LAYER QB ;
        RECT 61.2 0 66 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER JV ;
      RECT 0 0 80 60 ;
    LAYER YS ;
      RECT 0 0 80 60 ;
    LAYER JW ;
      RECT 0 0 80 60 ;
    LAYER QB ;
      RECT 0 0 80 60 ;
    LAYER QA ;
      RECT 0 0 80 60 ;
    LAYER JA ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_IO_SIG_H

MACRO RIIO_BUMP_RCUP100_DY
  CLASS COVER ;
  ORIGIN 30 30 ;
  FOREIGN RIIO_BUMP_RCUP100_DY -30 -30 ;
  SIZE 60 BY 60 ;
  SYMMETRY X Y R90 ;
  PIN DUMMY
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT -30 -13.713 30 13.713 ;
        RECT -25 -17.5 27.426 17.5 ;
        RECT -20 -22.5 22.426 22.5 ;
        RECT -15 -27.5 17.426 27.5 ;
        RECT -12.426 -30 12.426 30 ;
        RECT -15 -28.713 12.426 28.713 ;
        RECT -20 -24.926 17.426 24.926 ;
        RECT -25 -19.926 22.426 19.926 ;
        RECT -30 -14.926 27.426 14.926 ;
    END
  END DUMMY
  OBS
    LAYER LB ;
      RECT -12.426 -30 12.426 30 ;
      RECT -13.713 -29.357 12.426 29.357 ;
      RECT -13.713 -28.75 14.926 28.75 ;
      RECT -15 -28.713 14.926 28.713 ;
      RECT -15 -27.5 17.426 27.5 ;
      RECT -17.5 -26.176 17.426 26.176 ;
      RECT -20 -24.926 17.426 24.926 ;
      RECT -20 -23.75 19.926 23.75 ;
      RECT -20 -22.5 22.426 22.5 ;
      RECT -22.5 -21.176 22.426 21.176 ;
      RECT -25 -19.926 22.426 19.926 ;
      RECT -25 -18.75 24.926 18.75 ;
      RECT -25 -17.5 27.426 17.5 ;
      RECT -27.5 -16.176 27.426 16.176 ;
      RECT -30 -14.926 27.426 14.926 ;
      RECT -30 -14.357 28.713 14.357 ;
      RECT -30 -13.713 30 13.713 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  30 -14.379  28.047 -14.379  28.047 -16.332  26.094 -16.332  26.094 -18.284  24.142 -18.284  24.142 -20.237  22.189 -20.237  22.189 -22.19  20.236 -22.19  20.236 -24.142  18.284 -24.142  18.284 -26.095  16.331 -26.095  16.331 -28.048  14.378 -28.048  14.378 -30  -14.379 -30  -14.379 -28.047  -16.332 -28.047  -16.332 -26.094  -18.284 -26.094  -18.284 -24.142  -20.237 -24.142  -20.237 -22.189  -22.19 -22.189  -22.19 -20.236  -24.142 -20.236  -24.142 -18.284  -26.095 -18.284  -26.095 -16.331  -28.048 -16.331  -28.048 -14.378  -30 -14.378  -30 14.379  -28.047 14.379  -28.047 16.332  -26.094 16.332  -26.094 18.284  -24.142 18.284  -24.142 20.237  -22.189 20.237  -22.189 22.19  -20.236 22.19  -20.236 24.142  -18.284 24.142  -18.284 26.095  -16.331 26.095  -16.331 28.048  -14.378 28.048  -14.378 30  14.379 30  14.379 28.047  16.332 28.047  16.332 26.094  18.284 26.094  18.284 24.142  20.237 24.142  20.237 22.189  22.19 22.189  22.19 20.236  24.142 20.236  24.142 18.284  26.095 18.284  26.095 16.331  28.048 16.331  28.048 14.378  30 14.378 ;
  END
END RIIO_BUMP_RCUP100_DY

MACRO RIIO_BUMP_RCUP100_GND
  CLASS COVER ;
  ORIGIN 30 30 ;
  FOREIGN RIIO_BUMP_RCUP100_GND -30 -30 ;
  SIZE 60 BY 60 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 1.026 -13.713 30 13.713 ;
        RECT 1.026 -17.5 27.426 17.5 ;
        RECT 1.026 -22.5 22.426 22.5 ;
        RECT 1.026 -27.5 17.426 27.5 ;
        RECT -12.426 -8.974 12.426 30 ;
        RECT -12.426 -30 12.426 -11.026 ;
        RECT -30 -14.926 -1.026 14.926 ;
        RECT -15 -28.713 -1.026 28.713 ;
        RECT -20 -24.926 -1.026 24.926 ;
        RECT -25 -19.926 -1.026 19.926 ;
    END
  END VSS
  OBS
    LAYER LB ;
      RECT -12.426 -30 12.426 30 ;
      RECT -13.713 -29.357 12.426 29.357 ;
      RECT -13.713 -28.75 14.926 28.75 ;
      RECT -15 -28.713 14.926 28.713 ;
      RECT -15 -27.5 17.426 27.5 ;
      RECT -17.5 -26.176 17.426 26.176 ;
      RECT -20 -24.926 17.426 24.926 ;
      RECT -20 -23.75 19.926 23.75 ;
      RECT -20 -22.5 22.426 22.5 ;
      RECT -22.5 -21.176 22.426 21.176 ;
      RECT -25 -19.926 22.426 19.926 ;
      RECT -25 -18.75 24.926 18.75 ;
      RECT -25 -17.5 27.426 17.5 ;
      RECT -27.5 -16.176 27.426 16.176 ;
      RECT -30 -14.926 27.426 14.926 ;
      RECT -30 -14.357 28.713 14.357 ;
      RECT -30 -13.713 30 13.713 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  30 -14.379  28.047 -14.379  28.047 -16.332  26.094 -16.332  26.094 -18.284  24.142 -18.284  24.142 -20.237  22.189 -20.237  22.189 -22.19  20.236 -22.19  20.236 -24.142  18.284 -24.142  18.284 -26.095  16.331 -26.095  16.331 -28.048  14.378 -28.048  14.378 -30  -14.379 -30  -14.379 -28.047  -16.332 -28.047  -16.332 -26.094  -18.284 -26.094  -18.284 -24.142  -20.237 -24.142  -20.237 -22.189  -22.19 -22.189  -22.19 -20.236  -24.142 -20.236  -24.142 -18.284  -26.095 -18.284  -26.095 -16.331  -28.048 -16.331  -28.048 -14.378  -30 -14.378  -30 14.379  -28.047 14.379  -28.047 16.332  -26.094 16.332  -26.094 18.284  -24.142 18.284  -24.142 20.237  -22.189 20.237  -22.189 22.19  -20.236 22.19  -20.236 24.142  -18.284 24.142  -18.284 26.095  -16.331 26.095  -16.331 28.048  -14.378 28.048  -14.378 30  14.379 30  14.379 28.047  16.332 28.047  16.332 26.094  18.284 26.094  18.284 24.142  20.237 24.142  20.237 22.189  22.19 22.189  22.19 20.236  24.142 20.236  24.142 18.284  26.095 18.284  26.095 16.331  28.048 16.331  28.048 14.378  30 14.378 ;
  END
END RIIO_BUMP_RCUP100_GND

MACRO RIIO_BUMP_RCUP100_PWR
  CLASS COVER ;
  ORIGIN 30 30 ;
  FOREIGN RIIO_BUMP_RCUP100_PWR -30 -30 ;
  SIZE 60 BY 60 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 1.026 -13.713 30 13.713 ;
        RECT 1.026 -17.5 27.426 17.5 ;
        RECT 1.026 -22.5 22.426 22.5 ;
        RECT 1.026 -27.5 17.426 27.5 ;
        RECT -12.426 -8.974 12.426 30 ;
        RECT -12.426 -30 12.426 -11.026 ;
        RECT -30 -14.926 -1.026 14.926 ;
        RECT -15 -28.713 -1.026 28.713 ;
        RECT -20 -24.926 -1.026 24.926 ;
        RECT -25 -19.926 -1.026 19.926 ;
    END
  END VDD
  OBS
    LAYER LB ;
      RECT -12.426 -30 12.426 30 ;
      RECT -13.713 -29.357 12.426 29.357 ;
      RECT -13.713 -28.75 14.926 28.75 ;
      RECT -15 -28.713 14.926 28.713 ;
      RECT -15 -27.5 17.426 27.5 ;
      RECT -17.5 -26.176 17.426 26.176 ;
      RECT -20 -24.926 17.426 24.926 ;
      RECT -20 -23.75 19.926 23.75 ;
      RECT -20 -22.5 22.426 22.5 ;
      RECT -22.5 -21.176 22.426 21.176 ;
      RECT -25 -19.926 22.426 19.926 ;
      RECT -25 -18.75 24.926 18.75 ;
      RECT -25 -17.5 27.426 17.5 ;
      RECT -27.5 -16.176 27.426 16.176 ;
      RECT -30 -14.926 27.426 14.926 ;
      RECT -30 -14.357 28.713 14.357 ;
      RECT -30 -13.713 30 13.713 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  30 -14.379  28.047 -14.379  28.047 -16.332  26.094 -16.332  26.094 -18.284  24.142 -18.284  24.142 -20.237  22.189 -20.237  22.189 -22.19  20.236 -22.19  20.236 -24.142  18.284 -24.142  18.284 -26.095  16.331 -26.095  16.331 -28.048  14.378 -28.048  14.378 -30  -14.379 -30  -14.379 -28.047  -16.332 -28.047  -16.332 -26.094  -18.284 -26.094  -18.284 -24.142  -20.237 -24.142  -20.237 -22.189  -22.19 -22.189  -22.19 -20.236  -24.142 -20.236  -24.142 -18.284  -26.095 -18.284  -26.095 -16.331  -28.048 -16.331  -28.048 -14.378  -30 -14.378  -30 14.379  -28.047 14.379  -28.047 16.332  -26.094 16.332  -26.094 18.284  -24.142 18.284  -24.142 20.237  -22.189 20.237  -22.189 22.19  -20.236 22.19  -20.236 24.142  -18.284 24.142  -18.284 26.095  -16.331 26.095  -16.331 28.048  -14.378 28.048  -14.378 30  14.379 30  14.379 28.047  16.332 28.047  16.332 26.094  18.284 26.094  18.284 24.142  20.237 24.142  20.237 22.189  22.19 22.189  22.19 20.236  24.142 20.236  24.142 18.284  26.095 18.284  26.095 16.331  28.048 16.331  28.048 14.378  30 14.378 ;
  END
END RIIO_BUMP_RCUP100_PWR

MACRO RIIO_BUMP_RCUP100_SIG
  CLASS COVER ;
  ORIGIN 30 30 ;
  FOREIGN RIIO_BUMP_RCUP100_SIG -30 -30 ;
  SIZE 60 BY 60 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.210704 LAYER LB ;
    PORT
      LAYER LB ;
        RECT 1.026 -13.713 30 13.713 ;
        RECT 1.026 -17.5 27.426 17.5 ;
        RECT 1.026 -22.5 22.426 22.5 ;
        RECT 1.026 -27.5 17.426 27.5 ;
        RECT -12.426 -8.974 12.426 30 ;
        RECT -12.426 -30 12.426 -11.026 ;
        RECT -30 -14.926 -1.026 14.926 ;
        RECT -15 -28.713 -1.026 28.713 ;
        RECT -20 -24.926 -1.026 24.926 ;
        RECT -25 -19.926 -1.026 19.926 ;
    END
  END PAD
  OBS
    LAYER LB ;
      RECT -12.426 -30 12.426 30 ;
      RECT -13.713 -29.357 12.426 29.357 ;
      RECT -13.713 -28.75 14.926 28.75 ;
      RECT -15 -28.713 14.926 28.713 ;
      RECT -15 -27.5 17.426 27.5 ;
      RECT -17.5 -26.176 17.426 26.176 ;
      RECT -20 -24.926 17.426 24.926 ;
      RECT -20 -23.75 19.926 23.75 ;
      RECT -20 -22.5 22.426 22.5 ;
      RECT -22.5 -21.176 22.426 21.176 ;
      RECT -25 -19.926 22.426 19.926 ;
      RECT -25 -18.75 24.926 18.75 ;
      RECT -25 -17.5 27.426 17.5 ;
      RECT -27.5 -16.176 27.426 16.176 ;
      RECT -30 -14.926 27.426 14.926 ;
      RECT -30 -14.357 28.713 14.357 ;
      RECT -30 -13.713 30 13.713 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  30 -14.379  28.047 -14.379  28.047 -16.332  26.094 -16.332  26.094 -18.284  24.142 -18.284  24.142 -20.237  22.189 -20.237  22.189 -22.19  20.236 -22.19  20.236 -24.142  18.284 -24.142  18.284 -26.095  16.331 -26.095  16.331 -28.048  14.378 -28.048  14.378 -30  -14.379 -30  -14.379 -28.047  -16.332 -28.047  -16.332 -26.094  -18.284 -26.094  -18.284 -24.142  -20.237 -24.142  -20.237 -22.189  -22.19 -22.189  -22.19 -20.236  -24.142 -20.236  -24.142 -18.284  -26.095 -18.284  -26.095 -16.331  -28.048 -16.331  -28.048 -14.378  -30 -14.378  -30 14.379  -28.047 14.379  -28.047 16.332  -26.094 16.332  -26.094 18.284  -24.142 18.284  -24.142 20.237  -22.189 20.237  -22.189 22.19  -20.236 22.19  -20.236 24.142  -18.284 24.142  -18.284 26.095  -16.331 26.095  -16.331 28.048  -14.378 28.048  -14.378 30  14.379 30  14.379 28.047  16.332 28.047  16.332 26.094  18.284 26.094  18.284 24.142  20.237 24.142  20.237 22.189  22.19 22.189  22.19 20.236  24.142 20.236  24.142 18.284  26.095 18.284  26.095 16.331  28.048 16.331  28.048 14.378  30 14.378 ;
  END
END RIIO_BUMP_RCUP100_SIG

MACRO RIIO_BUMP_RCUP130_DY
  CLASS COVER ;
  ORIGIN 45 45 ;
  FOREIGN RIIO_BUMP_RCUP130_DY -45 -45 ;
  SIZE 90 BY 90 ;
  SYMMETRY X Y R90 ;
  PIN DUMMY
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT -45 -19.32 45 19.32 ;
        RECT -40 -22.5 43.639 22.5 ;
        RECT -35 -27.5 38.639 27.5 ;
        RECT -30 -32.5 33.639 32.5 ;
        RECT -25 -37.5 28.639 37.5 ;
        RECT -20 -42.5 23.639 42.5 ;
        RECT -18.639 -45 18.639 45 ;
        RECT -20 -44.32 18.639 44.32 ;
        RECT -25 -41.139 23.639 41.139 ;
        RECT -30 -36.139 28.639 36.139 ;
        RECT -35 -31.139 33.639 31.139 ;
        RECT -40 -26.139 38.639 26.139 ;
        RECT -45 -21.139 43.639 21.139 ;
    END
  END DUMMY
  OBS
    LAYER LB ;
      RECT -18.639 -45 18.639 45 ;
      RECT -19.319 -44.66 18.639 44.66 ;
      RECT -20 -44.32 18.639 44.32 ;
      RECT -20 -43.75 21.139 43.75 ;
      RECT -20 -42.5 23.639 42.5 ;
      RECT -22.5 -42.389 23.639 42.389 ;
      RECT -25 -41.139 23.639 41.139 ;
      RECT -25 -38.75 26.139 38.75 ;
      RECT -25 -37.5 28.639 37.5 ;
      RECT -27.5 -37.389 28.639 37.389 ;
      RECT -30 -36.139 28.639 36.139 ;
      RECT -30 -33.75 31.139 33.75 ;
      RECT -30 -32.5 33.639 32.5 ;
      RECT -32.5 -32.389 33.639 32.389 ;
      RECT -35 -31.139 33.639 31.139 ;
      RECT -35 -28.75 36.139 28.75 ;
      RECT -35 -27.5 38.639 27.5 ;
      RECT -37.5 -27.389 38.639 27.389 ;
      RECT -40 -26.139 38.639 26.139 ;
      RECT -40 -23.75 41.139 23.75 ;
      RECT -40 -22.5 43.639 22.5 ;
      RECT -42.5 -22.389 43.639 22.389 ;
      RECT -45 -21.139 43.639 21.139 ;
      RECT -45 -19.66 44.319 19.66 ;
      RECT -45 -19.32 45 19.32 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  45 -20.522  43.117 -20.522  43.117 -22.405  41.234 -22.405  41.234 -24.288  39.351 -24.288  39.351 -26.171  37.468 -26.171  37.468 -28.054  35.585 -28.054  35.585 -29.937  33.702 -29.937  33.702 -31.82  31.819 -31.82  31.819 -33.703  29.936 -33.703  29.936 -35.586  28.053 -35.586  28.053 -37.469  26.17 -37.469  26.17 -39.352  24.287 -39.352  24.287 -41.235  22.404 -41.235  22.404 -43.118  20.521 -43.118  20.521 -45  -20.522 -45  -20.522 -43.117  -22.405 -43.117  -22.405 -41.234  -24.288 -41.234  -24.288 -39.351  -26.171 -39.351  -26.171 -37.468  -28.054 -37.468  -28.054 -35.585  -29.937 -35.585  -29.937 -33.702  -31.82 -33.702  -31.82 -31.819  -33.703 -31.819  -33.703 -29.936  -35.586 -29.936  -35.586 -28.053  -37.469 -28.053  -37.469 -26.17  -39.352 -26.17  -39.352 -24.287  -41.235 -24.287  -41.235 -22.404  -43.118 -22.404  -43.118 -20.521  -45 -20.521  -45 20.522  -43.117 20.522  -43.117 22.405  -41.234 22.405  -41.234 24.288  -39.351 24.288  -39.351 26.171  -37.468 26.171  -37.468 28.054  -35.585 28.054  -35.585 29.937  -33.702 29.937  -33.702 31.82  -31.819 31.82  -31.819 33.703  -29.936 33.703  -29.936 35.586  -28.053 35.586  -28.053 37.469  -26.17 37.469  -26.17 39.352  -24.287 39.352  -24.287 41.235  -22.404 41.235  -22.404 43.118  -20.521 43.118  -20.521 45  20.522 45  20.522 43.117  22.405 43.117  22.405 41.234  24.288 41.234  24.288 39.351  26.171 39.351  26.171 37.468  28.054 37.468  28.054 35.585  29.937 35.585  29.937 33.702  31.82 33.702  31.82 31.819  33.703 31.819  33.703 29.936  35.586 29.936  35.586 28.053  37.469 28.053  37.469 26.17  39.352 26.17  39.352 24.287  41.235 24.287  41.235 22.404  43.118 22.404  43.118 20.521  45 20.521 ;
  END
END RIIO_BUMP_RCUP130_DY

MACRO RIIO_BUMP_RCUP130_GND
  CLASS COVER ;
  ORIGIN 45 45 ;
  FOREIGN RIIO_BUMP_RCUP130_GND -45 -45 ;
  SIZE 90 BY 90 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 1.026 -19.32 45 19.32 ;
        RECT 1.026 -22.5 43.639 22.5 ;
        RECT 1.026 -27.5 38.639 27.5 ;
        RECT 1.026 -32.5 33.639 32.5 ;
        RECT 1.026 -37.5 28.639 37.5 ;
        RECT 1.026 -42.5 23.639 42.5 ;
        RECT -18.639 -8.974 18.639 45 ;
        RECT -18.639 -45 18.639 -11.026 ;
        RECT -45 -21.139 -1.026 21.139 ;
        RECT -20 -44.32 -1.026 44.32 ;
        RECT -25 -41.139 -1.026 41.139 ;
        RECT -30 -36.139 -1.026 36.139 ;
        RECT -35 -31.139 -1.026 31.139 ;
        RECT -40 -26.139 -1.026 26.139 ;
    END
  END VSS
  OBS
    LAYER LB ;
      RECT -18.639 -45 18.639 45 ;
      RECT -19.319 -44.66 18.639 44.66 ;
      RECT -20 -44.32 18.639 44.32 ;
      RECT -20 -43.75 21.139 43.75 ;
      RECT -20 -42.5 23.639 42.5 ;
      RECT -22.5 -42.389 23.639 42.389 ;
      RECT -25 -41.139 23.639 41.139 ;
      RECT -25 -38.75 26.139 38.75 ;
      RECT -25 -37.5 28.639 37.5 ;
      RECT -27.5 -37.389 28.639 37.389 ;
      RECT -30 -36.139 28.639 36.139 ;
      RECT -30 -33.75 31.139 33.75 ;
      RECT -30 -32.5 33.639 32.5 ;
      RECT -32.5 -32.389 33.639 32.389 ;
      RECT -35 -31.139 33.639 31.139 ;
      RECT -35 -28.75 36.139 28.75 ;
      RECT -35 -27.5 38.639 27.5 ;
      RECT -37.5 -27.389 38.639 27.389 ;
      RECT -40 -26.139 38.639 26.139 ;
      RECT -40 -23.75 41.139 23.75 ;
      RECT -40 -22.5 43.639 22.5 ;
      RECT -42.5 -22.389 43.639 22.389 ;
      RECT -45 -21.139 43.639 21.139 ;
      RECT -45 -19.66 44.319 19.66 ;
      RECT -45 -19.32 45 19.32 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  45 -20.522  43.117 -20.522  43.117 -22.405  41.234 -22.405  41.234 -24.288  39.351 -24.288  39.351 -26.171  37.468 -26.171  37.468 -28.054  35.585 -28.054  35.585 -29.937  33.702 -29.937  33.702 -31.82  31.819 -31.82  31.819 -33.703  29.936 -33.703  29.936 -35.586  28.053 -35.586  28.053 -37.469  26.17 -37.469  26.17 -39.352  24.287 -39.352  24.287 -41.235  22.404 -41.235  22.404 -43.118  20.521 -43.118  20.521 -45  -20.522 -45  -20.522 -43.117  -22.405 -43.117  -22.405 -41.234  -24.288 -41.234  -24.288 -39.351  -26.171 -39.351  -26.171 -37.468  -28.054 -37.468  -28.054 -35.585  -29.937 -35.585  -29.937 -33.702  -31.82 -33.702  -31.82 -31.819  -33.703 -31.819  -33.703 -29.936  -35.586 -29.936  -35.586 -28.053  -37.469 -28.053  -37.469 -26.17  -39.352 -26.17  -39.352 -24.287  -41.235 -24.287  -41.235 -22.404  -43.118 -22.404  -43.118 -20.521  -45 -20.521  -45 20.522  -43.117 20.522  -43.117 22.405  -41.234 22.405  -41.234 24.288  -39.351 24.288  -39.351 26.171  -37.468 26.171  -37.468 28.054  -35.585 28.054  -35.585 29.937  -33.702 29.937  -33.702 31.82  -31.819 31.82  -31.819 33.703  -29.936 33.703  -29.936 35.586  -28.053 35.586  -28.053 37.469  -26.17 37.469  -26.17 39.352  -24.287 39.352  -24.287 41.235  -22.404 41.235  -22.404 43.118  -20.521 43.118  -20.521 45  20.522 45  20.522 43.117  22.405 43.117  22.405 41.234  24.288 41.234  24.288 39.351  26.171 39.351  26.171 37.468  28.054 37.468  28.054 35.585  29.937 35.585  29.937 33.702  31.82 33.702  31.82 31.819  33.703 31.819  33.703 29.936  35.586 29.936  35.586 28.053  37.469 28.053  37.469 26.17  39.352 26.17  39.352 24.287  41.235 24.287  41.235 22.404  43.118 22.404  43.118 20.521  45 20.521 ;
  END
END RIIO_BUMP_RCUP130_GND

MACRO RIIO_BUMP_RCUP130_PWR
  CLASS COVER ;
  ORIGIN 45 45 ;
  FOREIGN RIIO_BUMP_RCUP130_PWR -45 -45 ;
  SIZE 90 BY 90 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 1.026 -19.32 45 19.32 ;
        RECT 1.026 -22.5 43.639 22.5 ;
        RECT 1.026 -27.5 38.639 27.5 ;
        RECT 1.026 -32.5 33.639 32.5 ;
        RECT 1.026 -37.5 28.639 37.5 ;
        RECT 1.026 -42.5 23.639 42.5 ;
        RECT -18.639 -8.974 18.639 45 ;
        RECT -18.639 -45 18.639 -11.026 ;
        RECT -45 -21.139 -1.026 21.139 ;
        RECT -20 -44.32 -1.026 44.32 ;
        RECT -25 -41.139 -1.026 41.139 ;
        RECT -30 -36.139 -1.026 36.139 ;
        RECT -35 -31.139 -1.026 31.139 ;
        RECT -40 -26.139 -1.026 26.139 ;
    END
  END VDD
  OBS
    LAYER LB ;
      RECT -18.639 -45 18.639 45 ;
      RECT -19.319 -44.66 18.639 44.66 ;
      RECT -20 -44.32 18.639 44.32 ;
      RECT -20 -43.75 21.139 43.75 ;
      RECT -20 -42.5 23.639 42.5 ;
      RECT -22.5 -42.389 23.639 42.389 ;
      RECT -25 -41.139 23.639 41.139 ;
      RECT -25 -38.75 26.139 38.75 ;
      RECT -25 -37.5 28.639 37.5 ;
      RECT -27.5 -37.389 28.639 37.389 ;
      RECT -30 -36.139 28.639 36.139 ;
      RECT -30 -33.75 31.139 33.75 ;
      RECT -30 -32.5 33.639 32.5 ;
      RECT -32.5 -32.389 33.639 32.389 ;
      RECT -35 -31.139 33.639 31.139 ;
      RECT -35 -28.75 36.139 28.75 ;
      RECT -35 -27.5 38.639 27.5 ;
      RECT -37.5 -27.389 38.639 27.389 ;
      RECT -40 -26.139 38.639 26.139 ;
      RECT -40 -23.75 41.139 23.75 ;
      RECT -40 -22.5 43.639 22.5 ;
      RECT -42.5 -22.389 43.639 22.389 ;
      RECT -45 -21.139 43.639 21.139 ;
      RECT -45 -19.66 44.319 19.66 ;
      RECT -45 -19.32 45 19.32 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  45 -20.522  43.117 -20.522  43.117 -22.405  41.234 -22.405  41.234 -24.288  39.351 -24.288  39.351 -26.171  37.468 -26.171  37.468 -28.054  35.585 -28.054  35.585 -29.937  33.702 -29.937  33.702 -31.82  31.819 -31.82  31.819 -33.703  29.936 -33.703  29.936 -35.586  28.053 -35.586  28.053 -37.469  26.17 -37.469  26.17 -39.352  24.287 -39.352  24.287 -41.235  22.404 -41.235  22.404 -43.118  20.521 -43.118  20.521 -45  -20.522 -45  -20.522 -43.117  -22.405 -43.117  -22.405 -41.234  -24.288 -41.234  -24.288 -39.351  -26.171 -39.351  -26.171 -37.468  -28.054 -37.468  -28.054 -35.585  -29.937 -35.585  -29.937 -33.702  -31.82 -33.702  -31.82 -31.819  -33.703 -31.819  -33.703 -29.936  -35.586 -29.936  -35.586 -28.053  -37.469 -28.053  -37.469 -26.17  -39.352 -26.17  -39.352 -24.287  -41.235 -24.287  -41.235 -22.404  -43.118 -22.404  -43.118 -20.521  -45 -20.521  -45 20.522  -43.117 20.522  -43.117 22.405  -41.234 22.405  -41.234 24.288  -39.351 24.288  -39.351 26.171  -37.468 26.171  -37.468 28.054  -35.585 28.054  -35.585 29.937  -33.702 29.937  -33.702 31.82  -31.819 31.82  -31.819 33.703  -29.936 33.703  -29.936 35.586  -28.053 35.586  -28.053 37.469  -26.17 37.469  -26.17 39.352  -24.287 39.352  -24.287 41.235  -22.404 41.235  -22.404 43.118  -20.521 43.118  -20.521 45  20.522 45  20.522 43.117  22.405 43.117  22.405 41.234  24.288 41.234  24.288 39.351  26.171 39.351  26.171 37.468  28.054 37.468  28.054 35.585  29.937 35.585  29.937 33.702  31.82 33.702  31.82 31.819  33.703 31.819  33.703 29.936  35.586 29.936  35.586 28.053  37.469 28.053  37.469 26.17  39.352 26.17  39.352 24.287  41.235 24.287  41.235 22.404  43.118 22.404  43.118 20.521  45 20.521 ;
  END
END RIIO_BUMP_RCUP130_PWR

MACRO RIIO_BUMP_RCUP130_SIG
  CLASS COVER ;
  ORIGIN 45 45 ;
  FOREIGN RIIO_BUMP_RCUP130_SIG -45 -45 ;
  SIZE 90 BY 90 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.207982 LAYER LB ;
    PORT
      LAYER LB ;
        RECT 1.026 -19.32 45 19.32 ;
        RECT 1.026 -22.5 43.639 22.5 ;
        RECT 1.026 -27.5 38.639 27.5 ;
        RECT 1.026 -32.5 33.639 32.5 ;
        RECT 1.026 -37.5 28.639 37.5 ;
        RECT 1.026 -42.5 23.639 42.5 ;
        RECT -18.639 -8.974 18.639 45 ;
        RECT -18.639 -45 18.639 -11.026 ;
        RECT -45 -21.139 -1.026 21.139 ;
        RECT -20 -44.32 -1.026 44.32 ;
        RECT -25 -41.139 -1.026 41.139 ;
        RECT -30 -36.139 -1.026 36.139 ;
        RECT -35 -31.139 -1.026 31.139 ;
        RECT -40 -26.139 -1.026 26.139 ;
    END
  END PAD
  OBS
    LAYER LB ;
      RECT -18.639 -45 18.639 45 ;
      RECT -19.319 -44.66 18.639 44.66 ;
      RECT -20 -44.32 18.639 44.32 ;
      RECT -20 -43.75 21.139 43.75 ;
      RECT -20 -42.5 23.639 42.5 ;
      RECT -22.5 -42.389 23.639 42.389 ;
      RECT -25 -41.139 23.639 41.139 ;
      RECT -25 -38.75 26.139 38.75 ;
      RECT -25 -37.5 28.639 37.5 ;
      RECT -27.5 -37.389 28.639 37.389 ;
      RECT -30 -36.139 28.639 36.139 ;
      RECT -30 -33.75 31.139 33.75 ;
      RECT -30 -32.5 33.639 32.5 ;
      RECT -32.5 -32.389 33.639 32.389 ;
      RECT -35 -31.139 33.639 31.139 ;
      RECT -35 -28.75 36.139 28.75 ;
      RECT -35 -27.5 38.639 27.5 ;
      RECT -37.5 -27.389 38.639 27.389 ;
      RECT -40 -26.139 38.639 26.139 ;
      RECT -40 -23.75 41.139 23.75 ;
      RECT -40 -22.5 43.639 22.5 ;
      RECT -42.5 -22.389 43.639 22.389 ;
      RECT -45 -21.139 43.639 21.139 ;
      RECT -45 -19.66 44.319 19.66 ;
      RECT -45 -19.32 45 19.32 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  45 -20.522  43.117 -20.522  43.117 -22.405  41.234 -22.405  41.234 -24.288  39.351 -24.288  39.351 -26.171  37.468 -26.171  37.468 -28.054  35.585 -28.054  35.585 -29.937  33.702 -29.937  33.702 -31.82  31.819 -31.82  31.819 -33.703  29.936 -33.703  29.936 -35.586  28.053 -35.586  28.053 -37.469  26.17 -37.469  26.17 -39.352  24.287 -39.352  24.287 -41.235  22.404 -41.235  22.404 -43.118  20.521 -43.118  20.521 -45  -20.522 -45  -20.522 -43.117  -22.405 -43.117  -22.405 -41.234  -24.288 -41.234  -24.288 -39.351  -26.171 -39.351  -26.171 -37.468  -28.054 -37.468  -28.054 -35.585  -29.937 -35.585  -29.937 -33.702  -31.82 -33.702  -31.82 -31.819  -33.703 -31.819  -33.703 -29.936  -35.586 -29.936  -35.586 -28.053  -37.469 -28.053  -37.469 -26.17  -39.352 -26.17  -39.352 -24.287  -41.235 -24.287  -41.235 -22.404  -43.118 -22.404  -43.118 -20.521  -45 -20.521  -45 20.522  -43.117 20.522  -43.117 22.405  -41.234 22.405  -41.234 24.288  -39.351 24.288  -39.351 26.171  -37.468 26.171  -37.468 28.054  -35.585 28.054  -35.585 29.937  -33.702 29.937  -33.702 31.82  -31.819 31.82  -31.819 33.703  -29.936 33.703  -29.936 35.586  -28.053 35.586  -28.053 37.469  -26.17 37.469  -26.17 39.352  -24.287 39.352  -24.287 41.235  -22.404 41.235  -22.404 43.118  -20.521 43.118  -20.521 45  20.522 45  20.522 43.117  22.405 43.117  22.405 41.234  24.288 41.234  24.288 39.351  26.171 39.351  26.171 37.468  28.054 37.468  28.054 35.585  29.937 35.585  29.937 33.702  31.82 33.702  31.82 31.819  33.703 31.819  33.703 29.936  35.586 29.936  35.586 28.053  37.469 28.053  37.469 26.17  39.352 26.17  39.352 24.287  41.235 24.287  41.235 22.404  43.118 22.404  43.118 20.521  45 20.521 ;
  END
END RIIO_BUMP_RCUP130_SIG

MACRO RIIO_BUMP_SNAG140_DY
  CLASS COVER ;
  ORIGIN 35.5 35.5 ;
  FOREIGN RIIO_BUMP_SNAG140_DY -35.5 -35.5 ;
  SIZE 71 BY 71 ;
  SYMMETRY X Y R90 ;
  PIN DUMMY
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT -35.5 -15.103 35.5 15.103 ;
        RECT -30.5 -18 34.705 18 ;
        RECT -25.5 -23 29.705 23 ;
        RECT -20.5 -28 24.705 28 ;
        RECT -15.5 -33 19.705 33 ;
        RECT -14.705 -35.5 14.705 35.5 ;
        RECT -15.5 -35.103 14.705 35.103 ;
        RECT -20.5 -32.205 19.705 32.205 ;
        RECT -25.5 -27.205 24.705 27.205 ;
        RECT -30.5 -22.205 29.705 22.205 ;
        RECT -35.5 -17.205 34.705 17.205 ;
    END
  END DUMMY
  OBS
    LAYER LB ;
      RECT -14.705 -35.5 14.705 35.5 ;
      RECT -15.102 -35.302 14.705 35.302 ;
      RECT -15.5 -35.103 14.705 35.103 ;
      RECT -15.5 -34.25 17.205 34.25 ;
      RECT -18 -33.455 17.205 33.455 ;
      RECT -18 -33 19.705 33 ;
      RECT -20.5 -32.205 19.705 32.205 ;
      RECT -20.5 -29.25 22.205 29.25 ;
      RECT -23 -28.455 22.205 28.455 ;
      RECT -23 -28 24.705 28 ;
      RECT -25.5 -27.205 24.705 27.205 ;
      RECT -25.5 -24.25 27.205 24.25 ;
      RECT -28 -23.455 27.205 23.455 ;
      RECT -28 -23 29.705 23 ;
      RECT -30.5 -22.205 29.705 22.205 ;
      RECT -30.5 -19.25 32.205 19.25 ;
      RECT -33 -18.455 32.205 18.455 ;
      RECT -33 -18 34.705 18 ;
      RECT -35.5 -17.205 34.705 17.205 ;
      RECT -35.5 -15.302 35.102 15.302 ;
      RECT -35.5 -15.103 35.5 15.103 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  35.5 -16.596  33.609 -16.596  33.609 -18.486  31.719 -18.486  31.719 -20.377  29.828 -20.377  29.828 -22.267  27.938 -22.267  27.938 -24.158  26.047 -24.158  26.047 -26.048  24.157 -26.048  24.157 -27.939  22.266 -27.939  22.266 -29.829  20.376 -29.829  20.376 -31.72  18.485 -31.72  18.485 -33.61  16.595 -33.61  16.595 -35.5  -16.596 -35.5  -16.596 -33.609  -18.486 -33.609  -18.486 -31.719  -20.377 -31.719  -20.377 -29.828  -22.267 -29.828  -22.267 -27.938  -24.158 -27.938  -24.158 -26.047  -26.048 -26.047  -26.048 -24.157  -27.939 -24.157  -27.939 -22.266  -29.829 -22.266  -29.829 -20.376  -31.72 -20.376  -31.72 -18.485  -33.61 -18.485  -33.61 -16.595  -35.5 -16.595  -35.5 16.596  -33.609 16.596  -33.609 18.486  -31.719 18.486  -31.719 20.377  -29.828 20.377  -29.828 22.267  -27.938 22.267  -27.938 24.158  -26.047 24.158  -26.047 26.048  -24.157 26.048  -24.157 27.939  -22.266 27.939  -22.266 29.829  -20.376 29.829  -20.376 31.72  -18.485 31.72  -18.485 33.61  -16.595 33.61  -16.595 35.5  16.596 35.5  16.596 33.609  18.486 33.609  18.486 31.719  20.377 31.719  20.377 29.828  22.267 29.828  22.267 27.938  24.158 27.938  24.158 26.047  26.048 26.047  26.048 24.157  27.939 24.157  27.939 22.266  29.829 22.266  29.829 20.376  31.72 20.376  31.72 18.485  33.61 18.485  33.61 16.595  35.5 16.595 ;
  END
END RIIO_BUMP_SNAG140_DY

MACRO RIIO_BUMP_SNAG140_GND
  CLASS COVER ;
  ORIGIN 35.5 35.5 ;
  FOREIGN RIIO_BUMP_SNAG140_GND -35.5 -35.5 ;
  SIZE 71 BY 71 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 1.026 -15.102 35.5 15.103 ;
        RECT 1.026 -17.999 34.705 18 ;
        RECT 1.026 -22.999 29.705 23 ;
        RECT 1.026 -27.999 24.705 28 ;
        RECT 1.026 -32.999 19.705 33 ;
        RECT -14.705 -8.974 14.705 35.5 ;
        RECT 1.026 -35.499 14.705 35.5 ;
        RECT -14.705 -35.5 14.704 -11.026 ;
        RECT -35.5 -17.205 -1.026 17.205 ;
        RECT -15.5 -35.103 -1.026 35.103 ;
        RECT -20.5 -32.205 -1.026 32.205 ;
        RECT -25.5 -27.205 -1.026 27.205 ;
        RECT -30.5 -22.205 -1.026 22.205 ;
    END
  END VSS
  OBS
    LAYER LB ;
      RECT -14.705 -35.5 14.705 35.5 ;
      RECT -15.102 -35.302 14.705 35.302 ;
      RECT -15.5 -35.103 14.705 35.103 ;
      RECT -15.5 -34.25 17.205 34.25 ;
      RECT -18 -33.455 17.205 33.455 ;
      RECT -18 -32.999 19.705 33 ;
      RECT -20.5 -32.205 19.705 32.205 ;
      RECT -20.5 -29.25 22.205 29.25 ;
      RECT -23 -28.455 22.205 28.455 ;
      RECT -23 -27.999 24.705 28 ;
      RECT -25.5 -27.205 24.705 27.205 ;
      RECT -25.5 -24.25 27.205 24.25 ;
      RECT -28 -23.455 27.205 23.455 ;
      RECT -28 -22.999 29.705 23 ;
      RECT -30.5 -22.205 29.705 22.205 ;
      RECT -30.5 -19.25 32.205 19.25 ;
      RECT -33 -18.455 32.205 18.455 ;
      RECT -33 -17.999 34.705 18 ;
      RECT -35.5 -17.205 34.705 17.205 ;
      RECT -35.5 -15.302 35.102 15.302 ;
      RECT -35.5 -15.102 35.5 15.103 ;
      RECT -35.5 -15.103 35.103 15.103 ;
      RECT -33 -18 32.206 18 ;
      RECT -28 -23 27.206 23 ;
      RECT -23 -28 22.206 28 ;
      RECT -18 -33 17.206 33 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  35.5 -16.596  33.609 -16.596  33.609 -18.486  31.719 -18.486  31.719 -20.377  29.828 -20.377  29.828 -22.267  27.938 -22.267  27.938 -24.158  26.047 -24.158  26.047 -26.048  24.157 -26.048  24.157 -27.939  22.266 -27.939  22.266 -29.829  20.376 -29.829  20.376 -31.72  18.485 -31.72  18.485 -33.61  16.595 -33.61  16.595 -35.5  -16.596 -35.5  -16.596 -33.609  -18.486 -33.609  -18.486 -31.719  -20.377 -31.719  -20.377 -29.828  -22.267 -29.828  -22.267 -27.938  -24.158 -27.938  -24.158 -26.047  -26.048 -26.047  -26.048 -24.157  -27.939 -24.157  -27.939 -22.266  -29.829 -22.266  -29.829 -20.376  -31.72 -20.376  -31.72 -18.485  -33.61 -18.485  -33.61 -16.595  -35.5 -16.595  -35.5 16.596  -33.609 16.596  -33.609 18.486  -31.719 18.486  -31.719 20.377  -29.828 20.377  -29.828 22.267  -27.938 22.267  -27.938 24.158  -26.047 24.158  -26.047 26.048  -24.157 26.048  -24.157 27.939  -22.266 27.939  -22.266 29.829  -20.376 29.829  -20.376 31.72  -18.485 31.72  -18.485 33.61  -16.595 33.61  -16.595 35.5  16.596 35.5  16.596 33.609  18.486 33.609  18.486 31.719  20.377 31.719  20.377 29.828  22.267 29.828  22.267 27.938  24.158 27.938  24.158 26.047  26.048 26.047  26.048 24.157  27.939 24.157  27.939 22.266  29.829 22.266  29.829 20.376  31.72 20.376  31.72 18.485  33.61 18.485  33.61 16.595  35.5 16.595 ;
  END
END RIIO_BUMP_SNAG140_GND

MACRO RIIO_BUMP_SNAG140_PWR
  CLASS COVER ;
  ORIGIN 35.5 35.5 ;
  FOREIGN RIIO_BUMP_SNAG140_PWR -35.5 -35.5 ;
  SIZE 71 BY 71 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 1.026 -15.102 35.5 15.103 ;
        RECT 1.026 -17.999 34.705 18 ;
        RECT 1.026 -22.999 29.705 23 ;
        RECT 1.026 -27.999 24.705 28 ;
        RECT 1.026 -32.999 19.705 33 ;
        RECT -14.705 -8.974 14.705 35.5 ;
        RECT 1.026 -35.499 14.705 35.5 ;
        RECT -14.705 -35.5 14.704 -11.026 ;
        RECT -35.5 -17.205 -1.026 17.205 ;
        RECT -15.5 -35.103 -1.026 35.103 ;
        RECT -20.5 -32.205 -1.026 32.205 ;
        RECT -25.5 -27.205 -1.026 27.205 ;
        RECT -30.5 -22.205 -1.026 22.205 ;
    END
  END VDD
  OBS
    LAYER LB ;
      RECT -14.705 -35.5 14.705 35.5 ;
      RECT -15.102 -35.302 14.705 35.302 ;
      RECT -15.5 -35.103 14.705 35.103 ;
      RECT -15.5 -34.25 17.205 34.25 ;
      RECT -18 -33.455 17.205 33.455 ;
      RECT -18 -32.999 19.705 33 ;
      RECT -20.5 -32.205 19.705 32.205 ;
      RECT -20.5 -29.25 22.205 29.25 ;
      RECT -23 -28.455 22.205 28.455 ;
      RECT -23 -27.999 24.705 28 ;
      RECT -25.5 -27.205 24.705 27.205 ;
      RECT -25.5 -24.25 27.205 24.25 ;
      RECT -28 -23.455 27.205 23.455 ;
      RECT -28 -22.999 29.705 23 ;
      RECT -30.5 -22.205 29.705 22.205 ;
      RECT -30.5 -19.25 32.205 19.25 ;
      RECT -33 -18.455 32.205 18.455 ;
      RECT -33 -17.999 34.705 18 ;
      RECT -35.5 -17.205 34.705 17.205 ;
      RECT -35.5 -15.302 35.102 15.302 ;
      RECT -35.5 -15.102 35.5 15.103 ;
      RECT -35.5 -15.103 35.103 15.103 ;
      RECT -33 -18 32.206 18 ;
      RECT -28 -23 27.206 23 ;
      RECT -23 -28 22.206 28 ;
      RECT -18 -33 17.206 33 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  35.5 -16.596  33.609 -16.596  33.609 -18.486  31.719 -18.486  31.719 -20.377  29.828 -20.377  29.828 -22.267  27.938 -22.267  27.938 -24.158  26.047 -24.158  26.047 -26.048  24.157 -26.048  24.157 -27.939  22.266 -27.939  22.266 -29.829  20.376 -29.829  20.376 -31.72  18.485 -31.72  18.485 -33.61  16.595 -33.61  16.595 -35.5  -16.596 -35.5  -16.596 -33.609  -18.486 -33.609  -18.486 -31.719  -20.377 -31.719  -20.377 -29.828  -22.267 -29.828  -22.267 -27.938  -24.158 -27.938  -24.158 -26.047  -26.048 -26.047  -26.048 -24.157  -27.939 -24.157  -27.939 -22.266  -29.829 -22.266  -29.829 -20.376  -31.72 -20.376  -31.72 -18.485  -33.61 -18.485  -33.61 -16.595  -35.5 -16.595  -35.5 16.596  -33.609 16.596  -33.609 18.486  -31.719 18.486  -31.719 20.377  -29.828 20.377  -29.828 22.267  -27.938 22.267  -27.938 24.158  -26.047 24.158  -26.047 26.048  -24.157 26.048  -24.157 27.939  -22.266 27.939  -22.266 29.829  -20.376 29.829  -20.376 31.72  -18.485 31.72  -18.485 33.61  -16.595 33.61  -16.595 35.5  16.596 35.5  16.596 33.609  18.486 33.609  18.486 31.719  20.377 31.719  20.377 29.828  22.267 29.828  22.267 27.938  24.158 27.938  24.158 26.047  26.048 26.047  26.048 24.157  27.939 24.157  27.939 22.266  29.829 22.266  29.829 20.376  31.72 20.376  31.72 18.485  33.61 18.485  33.61 16.595  35.5 16.595 ;
  END
END RIIO_BUMP_SNAG140_PWR

MACRO RIIO_BUMP_SNAG140_SIG
  CLASS COVER ;
  ORIGIN 35.5 35.5 ;
  FOREIGN RIIO_BUMP_SNAG140_SIG -35.5 -35.5 ;
  SIZE 71 BY 71 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.22991 LAYER LB ;
    PORT
      LAYER LB ;
        RECT 1.026 -15.102 35.5 15.103 ;
        RECT 1.026 -17.999 34.705 18 ;
        RECT 1.026 -22.999 29.705 23 ;
        RECT 1.026 -27.999 24.705 28 ;
        RECT 1.026 -32.999 19.705 33 ;
        RECT -14.705 -8.974 14.705 35.5 ;
        RECT 1.026 -35.499 14.705 35.5 ;
        RECT -14.705 -35.5 14.704 -11.026 ;
        RECT -35.5 -17.205 -1.026 17.205 ;
        RECT -15.5 -35.103 -1.026 35.103 ;
        RECT -20.5 -32.205 -1.026 32.205 ;
        RECT -25.5 -27.205 -1.026 27.205 ;
        RECT -30.5 -22.205 -1.026 22.205 ;
    END
  END PAD
  OBS
    LAYER LB ;
      RECT -14.705 -35.5 14.705 35.5 ;
      RECT -15.102 -35.302 14.705 35.302 ;
      RECT -15.5 -35.103 14.705 35.103 ;
      RECT -15.5 -34.25 17.205 34.25 ;
      RECT -18 -33.455 17.205 33.455 ;
      RECT -18 -32.999 19.705 33 ;
      RECT -20.5 -32.205 19.705 32.205 ;
      RECT -20.5 -29.25 22.205 29.25 ;
      RECT -23 -28.455 22.205 28.455 ;
      RECT -23 -27.999 24.705 28 ;
      RECT -25.5 -27.205 24.705 27.205 ;
      RECT -25.5 -24.25 27.205 24.25 ;
      RECT -28 -23.455 27.205 23.455 ;
      RECT -28 -22.999 29.705 23 ;
      RECT -30.5 -22.205 29.705 22.205 ;
      RECT -30.5 -19.25 32.205 19.25 ;
      RECT -33 -18.455 32.205 18.455 ;
      RECT -33 -17.999 34.705 18 ;
      RECT -35.5 -17.205 34.705 17.205 ;
      RECT -35.5 -15.302 35.102 15.302 ;
      RECT -35.5 -15.102 35.5 15.103 ;
      RECT -35.5 -15.103 35.103 15.103 ;
      RECT -33 -18 32.206 18 ;
      RECT -28 -23 27.206 23 ;
      RECT -23 -28 22.206 28 ;
      RECT -18 -33 17.206 33 ;
    LAYER VV ;
      RECT -12.012 -29 12.012 29 ;
      RECT -14 -28.006 12.012 28.006 ;
      RECT -14 -26.5 17.012 26.5 ;
      RECT -19 -24.512 17.012 24.512 ;
      RECT -19 -21.5 22.012 21.5 ;
      RECT -24 -19.512 22.012 19.512 ;
      RECT -24 -16.5 27.012 16.5 ;
      RECT -29 -14.512 27.012 14.512 ;
      RECT -29 -13.006 29 13.006 ;
    LAYER OVERLAP ;
      POLYGON  35.5 -16.596  33.609 -16.596  33.609 -18.486  31.719 -18.486  31.719 -20.377  29.828 -20.377  29.828 -22.267  27.938 -22.267  27.938 -24.158  26.047 -24.158  26.047 -26.048  24.157 -26.048  24.157 -27.939  22.266 -27.939  22.266 -29.829  20.376 -29.829  20.376 -31.72  18.485 -31.72  18.485 -33.61  16.595 -33.61  16.595 -35.5  -16.596 -35.5  -16.596 -33.609  -18.486 -33.609  -18.486 -31.719  -20.377 -31.719  -20.377 -29.828  -22.267 -29.828  -22.267 -27.938  -24.158 -27.938  -24.158 -26.047  -26.048 -26.047  -26.048 -24.157  -27.939 -24.157  -27.939 -22.266  -29.829 -22.266  -29.829 -20.376  -31.72 -20.376  -31.72 -18.485  -33.61 -18.485  -33.61 -16.595  -35.5 -16.595  -35.5 16.596  -33.609 16.596  -33.609 18.486  -31.719 18.486  -31.719 20.377  -29.828 20.377  -29.828 22.267  -27.938 22.267  -27.938 24.158  -26.047 24.158  -26.047 26.048  -24.157 26.048  -24.157 27.939  -22.266 27.939  -22.266 29.829  -20.376 29.829  -20.376 31.72  -18.485 31.72  -18.485 33.61  -16.595 33.61  -16.595 35.5  16.596 35.5  16.596 33.609  18.486 33.609  18.486 31.719  20.377 31.719  20.377 29.828  22.267 29.828  22.267 27.938  24.158 27.938  24.158 26.047  26.048 26.047  26.048 24.157  27.939 24.157  27.939 22.266  29.829 22.266  29.829 20.376  31.72 20.376  31.72 18.485  33.61 18.485  33.61 16.595  35.5 16.595 ;
  END
END RIIO_BUMP_SNAG140_SIG

MACRO RIIO_BUMP_SNAG150_DY
  CLASS COVER ;
  ORIGIN 40.8 40.8 ;
  FOREIGN RIIO_BUMP_SNAG150_DY -40.8 -40.8 ;
  SIZE 81.6 BY 81.6 ;
  SYMMETRY X Y R90 ;
  PIN DUMMY
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT -40.8 -18.85 40.8 18.85 ;
        RECT -35.8 -23.3 36.9 23.3 ;
        RECT -30.8 -28.3 31.9 28.3 ;
        RECT -25.8 -33.3 26.9 33.3 ;
        RECT -20.8 -38.3 21.9 38.3 ;
        RECT -16.9 -40.8 16.9 40.8 ;
        RECT -20.8 -38.85 16.9 38.85 ;
        RECT -25.8 -34.4 21.9 34.4 ;
        RECT -30.8 -29.4 26.9 29.4 ;
        RECT -35.8 -24.4 31.9 24.4 ;
        RECT -40.8 -19.4 36.9 19.4 ;
    END
  END DUMMY
  OBS
    LAYER LB ;
      RECT -16.9 -40.8 16.9 40.8 ;
      RECT -18.85 -39.825 16.9 39.825 ;
      RECT -18.85 -39.55 19.4 39.55 ;
      RECT -20.8 -38.85 19.4 38.85 ;
      RECT -20.8 -38.3 21.9 38.3 ;
      RECT -23.3 -35.65 21.9 35.65 ;
      RECT -23.3 -34.55 24.4 34.55 ;
      RECT -25.8 -34.4 24.4 34.4 ;
      RECT -25.8 -33.3 26.9 33.3 ;
      RECT -28.3 -30.65 26.9 30.65 ;
      RECT -28.3 -29.55 29.4 29.55 ;
      RECT -30.8 -29.4 29.4 29.4 ;
      RECT -30.8 -28.3 31.9 28.3 ;
      RECT -33.3 -25.65 31.9 25.65 ;
      RECT -33.3 -24.55 34.4 24.55 ;
      RECT -35.8 -24.4 34.4 24.4 ;
      RECT -35.8 -23.3 36.9 23.3 ;
      RECT -38.3 -20.65 36.9 20.65 ;
      RECT -38.3 -19.825 38.85 19.825 ;
      RECT -40.8 -19.4 38.85 19.4 ;
      RECT -40.8 -18.85 40.8 18.85 ;
    LAYER VV ;
      RECT -15.533 -37.5 15.533 37.5 ;
      RECT -17.5 -36.517 15.533 36.517 ;
      RECT -17.5 -35 20.533 35 ;
      RECT -22.5 -33.033 20.533 33.033 ;
      RECT -22.5 -30 25.533 30 ;
      RECT -27.5 -28.033 25.533 28.033 ;
      RECT -27.5 -25 30.533 25 ;
      RECT -32.5 -23.033 30.533 23.033 ;
      RECT -32.5 -20 35.533 20 ;
      RECT -37.5 -18.033 35.533 18.033 ;
      RECT -37.5 -16.517 37.5 16.517 ;
    LAYER OVERLAP ;
      POLYGON  40.8 -18.892  38.808 -18.892  38.808 -20.884  36.816 -20.884  36.816 -22.875  34.825 -22.875  34.825 -24.867  32.833 -24.867  32.833 -26.859  30.841 -26.859  30.841 -28.85  28.85 -28.85  28.85 -30.842  26.858 -30.842  26.858 -32.834  24.866 -32.834  24.866 -34.825  22.875 -34.825  22.875 -36.817  20.883 -36.817  20.883 -38.809  18.891 -38.809  18.891 -40.8  -18.892 -40.8  -18.892 -38.808  -20.884 -38.808  -20.884 -36.816  -22.875 -36.816  -22.875 -34.825  -24.867 -34.825  -24.867 -32.833  -26.859 -32.833  -26.859 -30.841  -28.85 -30.841  -28.85 -28.85  -30.842 -28.85  -30.842 -26.858  -32.834 -26.858  -32.834 -24.866  -34.825 -24.866  -34.825 -22.875  -36.817 -22.875  -36.817 -20.883  -38.809 -20.883  -38.809 -18.891  -40.8 -18.891  -40.8 18.892  -38.808 18.892  -38.808 20.884  -36.816 20.884  -36.816 22.875  -34.825 22.875  -34.825 24.867  -32.833 24.867  -32.833 26.859  -30.841 26.859  -30.841 28.85  -28.85 28.85  -28.85 30.842  -26.858 30.842  -26.858 32.834  -24.866 32.834  -24.866 34.825  -22.875 34.825  -22.875 36.817  -20.883 36.817  -20.883 38.809  -18.891 38.809  -18.891 40.8  18.892 40.8  18.892 38.808  20.884 38.808  20.884 36.816  22.875 36.816  22.875 34.825  24.867 34.825  24.867 32.833  26.859 32.833  26.859 30.841  28.85 30.841  28.85 28.85  30.842 28.85  30.842 26.858  32.834 26.858  32.834 24.866  34.825 24.866  34.825 22.875  36.817 22.875  36.817 20.883  38.809 20.883  38.809 18.891  40.8 18.891 ;
  END
END RIIO_BUMP_SNAG150_DY

MACRO RIIO_BUMP_SNAG150_GND
  CLASS COVER ;
  ORIGIN 40.8 40.8 ;
  FOREIGN RIIO_BUMP_SNAG150_GND -40.8 -40.8 ;
  SIZE 81.6 BY 81.6 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 1.026 -18.85 40.8 18.85 ;
        RECT 1.026 -23.3 36.9 23.3 ;
        RECT 1.026 -28.3 31.9 28.3 ;
        RECT 1.026 -33.3 26.9 33.3 ;
        RECT 1.026 -38.3 21.9 38.3 ;
        RECT -16.9 -8.974 16.9 40.8 ;
        RECT -16.9 -40.8 16.9 -11.026 ;
        RECT -40.8 -19.4 -1.026 19.4 ;
        RECT -20.8 -38.85 -1.026 38.85 ;
        RECT -25.8 -34.4 -1.026 34.4 ;
        RECT -30.8 -29.4 -1.026 29.4 ;
        RECT -35.8 -24.4 -1.026 24.4 ;
    END
  END VSS
  OBS
    LAYER LB ;
      RECT -16.9 -40.8 16.9 40.8 ;
      RECT -18.85 -39.825 16.9 39.825 ;
      RECT -18.85 -39.55 19.4 39.55 ;
      RECT -20.8 -38.85 19.4 38.85 ;
      RECT -20.8 -38.3 21.9 38.3 ;
      RECT -23.3 -35.65 21.9 35.65 ;
      RECT -23.3 -34.55 24.4 34.55 ;
      RECT -25.8 -34.4 24.4 34.4 ;
      RECT -25.8 -33.3 26.9 33.3 ;
      RECT -28.3 -30.65 26.9 30.65 ;
      RECT -28.3 -29.55 29.4 29.55 ;
      RECT -30.8 -29.4 29.4 29.4 ;
      RECT -30.8 -28.3 31.9 28.3 ;
      RECT -33.3 -25.65 31.9 25.65 ;
      RECT -33.3 -24.55 34.4 24.55 ;
      RECT -35.8 -24.4 34.4 24.4 ;
      RECT -35.8 -23.3 36.9 23.3 ;
      RECT -38.3 -20.65 36.9 20.65 ;
      RECT -38.3 -19.825 38.85 19.825 ;
      RECT -40.8 -19.4 38.85 19.4 ;
      RECT -40.8 -18.85 40.8 18.85 ;
    LAYER VV ;
      RECT -15.533 -37.5 15.533 37.5 ;
      RECT -17.5 -36.517 15.533 36.517 ;
      RECT -17.5 -35 20.533 35 ;
      RECT -22.5 -33.033 20.533 33.033 ;
      RECT -22.5 -30 25.533 30 ;
      RECT -27.5 -28.033 25.533 28.033 ;
      RECT -27.5 -25 30.533 25 ;
      RECT -32.5 -23.033 30.533 23.033 ;
      RECT -32.5 -20 35.533 20 ;
      RECT -37.5 -18.033 35.533 18.033 ;
      RECT -37.5 -16.517 37.5 16.517 ;
    LAYER OVERLAP ;
      POLYGON  40.8 -18.892  38.808 -18.892  38.808 -20.884  36.816 -20.884  36.816 -22.875  34.825 -22.875  34.825 -24.867  32.833 -24.867  32.833 -26.859  30.841 -26.859  30.841 -28.85  28.85 -28.85  28.85 -30.842  26.858 -30.842  26.858 -32.834  24.866 -32.834  24.866 -34.825  22.875 -34.825  22.875 -36.817  20.883 -36.817  20.883 -38.809  18.891 -38.809  18.891 -40.8  -18.892 -40.8  -18.892 -38.808  -20.884 -38.808  -20.884 -36.816  -22.875 -36.816  -22.875 -34.825  -24.867 -34.825  -24.867 -32.833  -26.859 -32.833  -26.859 -30.841  -28.85 -30.841  -28.85 -28.85  -30.842 -28.85  -30.842 -26.858  -32.834 -26.858  -32.834 -24.866  -34.825 -24.866  -34.825 -22.875  -36.817 -22.875  -36.817 -20.883  -38.809 -20.883  -38.809 -18.891  -40.8 -18.891  -40.8 18.892  -38.808 18.892  -38.808 20.884  -36.816 20.884  -36.816 22.875  -34.825 22.875  -34.825 24.867  -32.833 24.867  -32.833 26.859  -30.841 26.859  -30.841 28.85  -28.85 28.85  -28.85 30.842  -26.858 30.842  -26.858 32.834  -24.866 32.834  -24.866 34.825  -22.875 34.825  -22.875 36.817  -20.883 36.817  -20.883 38.809  -18.891 38.809  -18.891 40.8  18.892 40.8  18.892 38.808  20.884 38.808  20.884 36.816  22.875 36.816  22.875 34.825  24.867 34.825  24.867 32.833  26.859 32.833  26.859 30.841  28.85 30.841  28.85 28.85  30.842 28.85  30.842 26.858  32.834 26.858  32.834 24.866  34.825 24.866  34.825 22.875  36.817 22.875  36.817 20.883  38.809 20.883  38.809 18.891  40.8 18.891 ;
  END
END RIIO_BUMP_SNAG150_GND

MACRO RIIO_BUMP_SNAG150_PWR
  CLASS COVER ;
  ORIGIN 40.8 40.8 ;
  FOREIGN RIIO_BUMP_SNAG150_PWR -40.8 -40.8 ;
  SIZE 81.6 BY 81.6 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 1.026 -18.85 40.8 18.85 ;
        RECT 1.026 -23.3 36.9 23.3 ;
        RECT 1.026 -28.3 31.9 28.3 ;
        RECT 1.026 -33.3 26.9 33.3 ;
        RECT 1.026 -38.3 21.9 38.3 ;
        RECT -16.9 -8.974 16.9 40.8 ;
        RECT -16.9 -40.8 16.9 -11.026 ;
        RECT -40.8 -19.4 -1.026 19.4 ;
        RECT -20.8 -38.85 -1.026 38.85 ;
        RECT -25.8 -34.4 -1.026 34.4 ;
        RECT -30.8 -29.4 -1.026 29.4 ;
        RECT -35.8 -24.4 -1.026 24.4 ;
    END
  END VDD
  OBS
    LAYER LB ;
      RECT -16.9 -40.8 16.9 40.8 ;
      RECT -18.85 -39.825 16.9 39.825 ;
      RECT -18.85 -39.55 19.4 39.55 ;
      RECT -20.8 -38.85 19.4 38.85 ;
      RECT -20.8 -38.3 21.9 38.3 ;
      RECT -23.3 -35.65 21.9 35.65 ;
      RECT -23.3 -34.55 24.4 34.55 ;
      RECT -25.8 -34.4 24.4 34.4 ;
      RECT -25.8 -33.3 26.9 33.3 ;
      RECT -28.3 -30.65 26.9 30.65 ;
      RECT -28.3 -29.55 29.4 29.55 ;
      RECT -30.8 -29.4 29.4 29.4 ;
      RECT -30.8 -28.3 31.9 28.3 ;
      RECT -33.3 -25.65 31.9 25.65 ;
      RECT -33.3 -24.55 34.4 24.55 ;
      RECT -35.8 -24.4 34.4 24.4 ;
      RECT -35.8 -23.3 36.9 23.3 ;
      RECT -38.3 -20.65 36.9 20.65 ;
      RECT -38.3 -19.825 38.85 19.825 ;
      RECT -40.8 -19.4 38.85 19.4 ;
      RECT -40.8 -18.85 40.8 18.85 ;
    LAYER VV ;
      RECT -15.533 -37.5 15.533 37.5 ;
      RECT -17.5 -36.517 15.533 36.517 ;
      RECT -17.5 -35 20.533 35 ;
      RECT -22.5 -33.033 20.533 33.033 ;
      RECT -22.5 -30 25.533 30 ;
      RECT -27.5 -28.033 25.533 28.033 ;
      RECT -27.5 -25 30.533 25 ;
      RECT -32.5 -23.033 30.533 23.033 ;
      RECT -32.5 -20 35.533 20 ;
      RECT -37.5 -18.033 35.533 18.033 ;
      RECT -37.5 -16.517 37.5 16.517 ;
    LAYER OVERLAP ;
      POLYGON  40.8 -18.892  38.808 -18.892  38.808 -20.884  36.816 -20.884  36.816 -22.875  34.825 -22.875  34.825 -24.867  32.833 -24.867  32.833 -26.859  30.841 -26.859  30.841 -28.85  28.85 -28.85  28.85 -30.842  26.858 -30.842  26.858 -32.834  24.866 -32.834  24.866 -34.825  22.875 -34.825  22.875 -36.817  20.883 -36.817  20.883 -38.809  18.891 -38.809  18.891 -40.8  -18.892 -40.8  -18.892 -38.808  -20.884 -38.808  -20.884 -36.816  -22.875 -36.816  -22.875 -34.825  -24.867 -34.825  -24.867 -32.833  -26.859 -32.833  -26.859 -30.841  -28.85 -30.841  -28.85 -28.85  -30.842 -28.85  -30.842 -26.858  -32.834 -26.858  -32.834 -24.866  -34.825 -24.866  -34.825 -22.875  -36.817 -22.875  -36.817 -20.883  -38.809 -20.883  -38.809 -18.891  -40.8 -18.891  -40.8 18.892  -38.808 18.892  -38.808 20.884  -36.816 20.884  -36.816 22.875  -34.825 22.875  -34.825 24.867  -32.833 24.867  -32.833 26.859  -30.841 26.859  -30.841 28.85  -28.85 28.85  -28.85 30.842  -26.858 30.842  -26.858 32.834  -24.866 32.834  -24.866 34.825  -22.875 34.825  -22.875 36.817  -20.883 36.817  -20.883 38.809  -18.891 38.809  -18.891 40.8  18.892 40.8  18.892 38.808  20.884 38.808  20.884 36.816  22.875 36.816  22.875 34.825  24.867 34.825  24.867 32.833  26.859 32.833  26.859 30.841  28.85 30.841  28.85 28.85  30.842 28.85  30.842 26.858  32.834 26.858  32.834 24.866  34.825 24.866  34.825 22.875  36.817 22.875  36.817 20.883  38.809 20.883  38.809 18.891  40.8 18.891 ;
  END
END RIIO_BUMP_SNAG150_PWR

MACRO RIIO_BUMP_SNAG150_SIG
  CLASS COVER ;
  ORIGIN 40.8 40.8 ;
  FOREIGN RIIO_BUMP_SNAG150_SIG -40.8 -40.8 ;
  SIZE 81.6 BY 81.6 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.210704 LAYER LB ;
    PORT
      LAYER LB ;
        RECT 1.026 -18.85 40.8 18.85 ;
        RECT 1.026 -23.3 36.9 23.3 ;
        RECT 1.026 -28.3 31.9 28.3 ;
        RECT 1.026 -33.3 26.9 33.3 ;
        RECT 1.026 -38.3 21.9 38.3 ;
        RECT -16.9 -8.974 16.9 40.8 ;
        RECT -16.9 -40.8 16.9 -11.026 ;
        RECT -40.8 -19.4 -1.026 19.4 ;
        RECT -20.8 -38.85 -1.026 38.85 ;
        RECT -25.8 -34.4 -1.026 34.4 ;
        RECT -30.8 -29.4 -1.026 29.4 ;
        RECT -35.8 -24.4 -1.026 24.4 ;
    END
  END PAD
  OBS
    LAYER LB ;
      RECT -16.9 -40.8 16.9 40.8 ;
      RECT -18.85 -39.825 16.9 39.825 ;
      RECT -18.85 -39.55 19.4 39.55 ;
      RECT -20.8 -38.85 19.4 38.85 ;
      RECT -20.8 -38.3 21.9 38.3 ;
      RECT -23.3 -35.65 21.9 35.65 ;
      RECT -23.3 -34.55 24.4 34.55 ;
      RECT -25.8 -34.4 24.4 34.4 ;
      RECT -25.8 -33.3 26.9 33.3 ;
      RECT -28.3 -30.65 26.9 30.65 ;
      RECT -28.3 -29.55 29.4 29.55 ;
      RECT -30.8 -29.4 29.4 29.4 ;
      RECT -30.8 -28.3 31.9 28.3 ;
      RECT -33.3 -25.65 31.9 25.65 ;
      RECT -33.3 -24.55 34.4 24.55 ;
      RECT -35.8 -24.4 34.4 24.4 ;
      RECT -35.8 -23.3 36.9 23.3 ;
      RECT -38.3 -20.65 36.9 20.65 ;
      RECT -38.3 -19.825 38.85 19.825 ;
      RECT -40.8 -19.4 38.85 19.4 ;
      RECT -40.8 -18.85 40.8 18.85 ;
    LAYER VV ;
      RECT -15.533 -37.5 15.533 37.5 ;
      RECT -17.5 -36.517 15.533 36.517 ;
      RECT -17.5 -35 20.533 35 ;
      RECT -22.5 -33.033 20.533 33.033 ;
      RECT -22.5 -30 25.533 30 ;
      RECT -27.5 -28.033 25.533 28.033 ;
      RECT -27.5 -25 30.533 25 ;
      RECT -32.5 -23.033 30.533 23.033 ;
      RECT -32.5 -20 35.533 20 ;
      RECT -37.5 -18.033 35.533 18.033 ;
      RECT -37.5 -16.517 37.5 16.517 ;
    LAYER OVERLAP ;
      POLYGON  40.8 -18.892  38.808 -18.892  38.808 -20.884  36.816 -20.884  36.816 -22.875  34.825 -22.875  34.825 -24.867  32.833 -24.867  32.833 -26.859  30.841 -26.859  30.841 -28.85  28.85 -28.85  28.85 -30.842  26.858 -30.842  26.858 -32.834  24.866 -32.834  24.866 -34.825  22.875 -34.825  22.875 -36.817  20.883 -36.817  20.883 -38.809  18.891 -38.809  18.891 -40.8  -18.892 -40.8  -18.892 -38.808  -20.884 -38.808  -20.884 -36.816  -22.875 -36.816  -22.875 -34.825  -24.867 -34.825  -24.867 -32.833  -26.859 -32.833  -26.859 -30.841  -28.85 -30.841  -28.85 -28.85  -30.842 -28.85  -30.842 -26.858  -32.834 -26.858  -32.834 -24.866  -34.825 -24.866  -34.825 -22.875  -36.817 -22.875  -36.817 -20.883  -38.809 -20.883  -38.809 -18.891  -40.8 -18.891  -40.8 18.892  -38.808 18.892  -38.808 20.884  -36.816 20.884  -36.816 22.875  -34.825 22.875  -34.825 24.867  -32.833 24.867  -32.833 26.859  -30.841 26.859  -30.841 28.85  -28.85 28.85  -28.85 30.842  -26.858 30.842  -26.858 32.834  -24.866 32.834  -24.866 34.825  -22.875 34.825  -22.875 36.817  -20.883 36.817  -20.883 38.809  -18.891 38.809  -18.891 40.8  18.892 40.8  18.892 38.808  20.884 38.808  20.884 36.816  22.875 36.816  22.875 34.825  24.867 34.825  24.867 32.833  26.859 32.833  26.859 30.841  28.85 30.841  28.85 28.85  30.842 28.85  30.842 26.858  32.834 26.858  32.834 24.866  34.825 24.866  34.825 22.875  36.817 22.875  36.817 20.883  38.809 20.883  38.809 18.891  40.8 18.891 ;
  END
END RIIO_BUMP_SNAG150_SIG

MACRO RIIO_BUMP_SNAG180_DY
  CLASS COVER ;
  ORIGIN 48 48 ;
  FOREIGN RIIO_BUMP_SNAG180_DY -48 -48 ;
  SIZE 96 BY 96 ;
  SYMMETRY X Y R90 ;
  PIN DUMMY
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT -48 -21.441 48 21.441 ;
        RECT -43 -25.5 44.882 25.5 ;
        RECT -38 -30.5 39.882 30.5 ;
        RECT -33 -35.5 34.882 35.5 ;
        RECT -28 -40.5 29.882 40.5 ;
        RECT -23 -45.5 24.882 45.5 ;
        RECT -19.882 -48 19.882 48 ;
        RECT -23 -46.441 19.882 46.441 ;
        RECT -28 -42.382 24.882 42.382 ;
        RECT -33 -37.382 29.882 37.382 ;
        RECT -38 -32.382 34.882 32.382 ;
        RECT -43 -27.382 39.882 27.382 ;
        RECT -48 -22.382 44.882 22.382 ;
    END
  END DUMMY
  OBS
    LAYER LB ;
      RECT -19.882 -48 19.882 48 ;
      RECT -21.441 -47.221 19.882 47.221 ;
      RECT -21.441 -46.75 22.382 46.75 ;
      RECT -23 -46.441 22.382 46.441 ;
      RECT -23 -45.5 24.882 45.5 ;
      RECT -25.5 -43.632 24.882 43.632 ;
      RECT -28 -42.382 24.882 42.382 ;
      RECT -28 -41.75 27.382 41.75 ;
      RECT -28 -40.5 29.882 40.5 ;
      RECT -30.5 -38.632 29.882 38.632 ;
      RECT -33 -37.382 29.882 37.382 ;
      RECT -33 -36.75 32.382 36.75 ;
      RECT -33 -35.5 34.882 35.5 ;
      RECT -35.5 -33.632 34.882 33.632 ;
      RECT -38 -32.382 34.882 32.382 ;
      RECT -38 -31.75 37.382 31.75 ;
      RECT -38 -30.5 39.882 30.5 ;
      RECT -40.5 -28.632 39.882 28.632 ;
      RECT -43 -27.382 39.882 27.382 ;
      RECT -43 -26.75 42.382 26.75 ;
      RECT -43 -25.5 44.882 25.5 ;
      RECT -45.5 -23.632 44.882 23.632 ;
      RECT -48 -22.382 44.882 22.382 ;
      RECT -48 -22.221 46.441 22.221 ;
      RECT -48 -21.441 48 21.441 ;
    LAYER VV ;
      RECT -19.261 -46.5 19.261 46.5 ;
      RECT -21.5 -45.381 19.261 45.381 ;
      RECT -21.5 -44 24.261 44 ;
      RECT -26.5 -41.761 24.261 41.761 ;
      RECT -26.5 -39 29.261 39 ;
      RECT -31.5 -36.761 29.261 36.761 ;
      RECT -31.5 -34 34.261 34 ;
      RECT -36.5 -31.761 34.261 31.761 ;
      RECT -36.5 -29 39.261 29 ;
      RECT -41.5 -26.761 39.261 26.761 ;
      RECT -41.5 -24 44.261 24 ;
      RECT -46.5 -21.761 44.261 21.761 ;
      RECT -46.5 -20.381 46.5 20.381 ;
    LAYER OVERLAP ;
      POLYGON  48 -21.757  46.125 -21.757  46.125 -23.632  44.25 -23.632  44.25 -25.506  42.376 -25.506  42.376 -27.381  40.501 -27.381  40.501 -29.255  38.627 -29.255  38.627 -31.13  36.752 -31.13  36.752 -33.004  34.878 -33.004  34.878 -34.879  33.003 -34.879  33.003 -36.753  31.129 -36.753  31.129 -38.628  29.254 -38.628  29.254 -40.502  27.38 -40.502  27.38 -42.377  25.505 -42.377  25.505 -44.251  23.631 -44.251  23.631 -46.126  21.756 -46.126  21.756 -48  -21.757 -48  -21.757 -46.125  -23.632 -46.125  -23.632 -44.25  -25.506 -44.25  -25.506 -42.376  -27.381 -42.376  -27.381 -40.501  -29.255 -40.501  -29.255 -38.627  -31.13 -38.627  -31.13 -36.752  -33.004 -36.752  -33.004 -34.878  -34.879 -34.878  -34.879 -33.003  -36.753 -33.003  -36.753 -31.129  -38.628 -31.129  -38.628 -29.254  -40.502 -29.254  -40.502 -27.38  -42.377 -27.38  -42.377 -25.505  -44.251 -25.505  -44.251 -23.631  -46.126 -23.631  -46.126 -21.756  -48 -21.756  -48 21.757  -46.125 21.757  -46.125 23.632  -44.25 23.632  -44.25 25.506  -42.376 25.506  -42.376 27.381  -40.501 27.381  -40.501 29.255  -38.627 29.255  -38.627 31.13  -36.752 31.13  -36.752 33.004  -34.878 33.004  -34.878 34.879  -33.003 34.879  -33.003 36.753  -31.129 36.753  -31.129 38.628  -29.254 38.628  -29.254 40.502  -27.38 40.502  -27.38 42.377  -25.505 42.377  -25.505 44.251  -23.631 44.251  -23.631 46.126  -21.756 46.126  -21.756 48  21.757 48  21.757 46.125  23.632 46.125  23.632 44.25  25.506 44.25  25.506 42.376  27.381 42.376  27.381 40.501  29.255 40.501  29.255 38.627  31.13 38.627  31.13 36.752  33.004 36.752  33.004 34.878  34.879 34.878  34.879 33.003  36.753 33.003  36.753 31.129  38.628 31.129  38.628 29.254  40.502 29.254  40.502 27.38  42.377 27.38  42.377 25.505  44.251 25.505  44.251 23.631  46.126 23.631  46.126 21.756  48 21.756 ;
  END
END RIIO_BUMP_SNAG180_DY

MACRO RIIO_BUMP_SNAG180_GND
  CLASS COVER ;
  ORIGIN 48 48 ;
  FOREIGN RIIO_BUMP_SNAG180_GND -48 -48 ;
  SIZE 96 BY 96 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 1.026 -21.441 48 21.441 ;
        RECT 1.026 -25.5 44.882 25.5 ;
        RECT 1.026 -30.5 39.882 30.5 ;
        RECT 1.026 -35.5 34.882 35.5 ;
        RECT 1.026 -40.5 29.882 40.5 ;
        RECT 1.026 -45.5 24.882 45.5 ;
        RECT -19.882 -8.974 19.882 48 ;
        RECT -19.882 -48 19.882 -11.026 ;
        RECT -48 -22.382 -1.026 22.382 ;
        RECT -23 -46.441 -1.026 46.441 ;
        RECT -28 -42.382 -1.026 42.382 ;
        RECT -33 -37.382 -1.026 37.382 ;
        RECT -38 -32.382 -1.026 32.382 ;
        RECT -43 -27.382 -1.026 27.382 ;
    END
  END VSS
  OBS
    LAYER LB ;
      RECT -19.882 -48 19.882 48 ;
      RECT -21.441 -47.221 19.882 47.221 ;
      RECT -21.441 -46.75 22.382 46.75 ;
      RECT -23 -46.441 22.382 46.441 ;
      RECT -23 -45.5 24.882 45.5 ;
      RECT -25.5 -43.632 24.882 43.632 ;
      RECT -28 -42.382 24.882 42.382 ;
      RECT -28 -41.75 27.382 41.75 ;
      RECT -28 -40.5 29.882 40.5 ;
      RECT -30.5 -38.632 29.882 38.632 ;
      RECT -33 -37.382 29.882 37.382 ;
      RECT -33 -36.75 32.382 36.75 ;
      RECT -33 -35.5 34.882 35.5 ;
      RECT -35.5 -33.632 34.882 33.632 ;
      RECT -38 -32.382 34.882 32.382 ;
      RECT -38 -31.75 37.382 31.75 ;
      RECT -38 -30.5 39.882 30.5 ;
      RECT -40.5 -28.632 39.882 28.632 ;
      RECT -43 -27.382 39.882 27.382 ;
      RECT -43 -26.75 42.382 26.75 ;
      RECT -43 -25.5 44.882 25.5 ;
      RECT -45.5 -23.632 44.882 23.632 ;
      RECT -48 -22.382 44.882 22.382 ;
      RECT -48 -22.221 46.441 22.221 ;
      RECT -48 -21.441 48 21.441 ;
    LAYER VV ;
      RECT -19.261 -46.5 19.261 46.5 ;
      RECT -21.5 -45.381 19.261 45.381 ;
      RECT -21.5 -44 24.261 44 ;
      RECT -26.5 -41.761 24.261 41.761 ;
      RECT -26.5 -39 29.261 39 ;
      RECT -31.5 -36.761 29.261 36.761 ;
      RECT -31.5 -34 34.261 34 ;
      RECT -36.5 -31.761 34.261 31.761 ;
      RECT -36.5 -29 39.261 29 ;
      RECT -41.5 -26.761 39.261 26.761 ;
      RECT -41.5 -24 44.261 24 ;
      RECT -46.5 -21.761 44.261 21.761 ;
      RECT -46.5 -20.381 46.5 20.381 ;
    LAYER OVERLAP ;
      POLYGON  48 -21.757  46.125 -21.757  46.125 -23.632  44.25 -23.632  44.25 -25.506  42.376 -25.506  42.376 -27.381  40.501 -27.381  40.501 -29.255  38.627 -29.255  38.627 -31.13  36.752 -31.13  36.752 -33.004  34.878 -33.004  34.878 -34.879  33.003 -34.879  33.003 -36.753  31.129 -36.753  31.129 -38.628  29.254 -38.628  29.254 -40.502  27.38 -40.502  27.38 -42.377  25.505 -42.377  25.505 -44.251  23.631 -44.251  23.631 -46.126  21.756 -46.126  21.756 -48  -21.757 -48  -21.757 -46.125  -23.632 -46.125  -23.632 -44.25  -25.506 -44.25  -25.506 -42.376  -27.381 -42.376  -27.381 -40.501  -29.255 -40.501  -29.255 -38.627  -31.13 -38.627  -31.13 -36.752  -33.004 -36.752  -33.004 -34.878  -34.879 -34.878  -34.879 -33.003  -36.753 -33.003  -36.753 -31.129  -38.628 -31.129  -38.628 -29.254  -40.502 -29.254  -40.502 -27.38  -42.377 -27.38  -42.377 -25.505  -44.251 -25.505  -44.251 -23.631  -46.126 -23.631  -46.126 -21.756  -48 -21.756  -48 21.757  -46.125 21.757  -46.125 23.632  -44.25 23.632  -44.25 25.506  -42.376 25.506  -42.376 27.381  -40.501 27.381  -40.501 29.255  -38.627 29.255  -38.627 31.13  -36.752 31.13  -36.752 33.004  -34.878 33.004  -34.878 34.879  -33.003 34.879  -33.003 36.753  -31.129 36.753  -31.129 38.628  -29.254 38.628  -29.254 40.502  -27.38 40.502  -27.38 42.377  -25.505 42.377  -25.505 44.251  -23.631 44.251  -23.631 46.126  -21.756 46.126  -21.756 48  21.757 48  21.757 46.125  23.632 46.125  23.632 44.25  25.506 44.25  25.506 42.376  27.381 42.376  27.381 40.501  29.255 40.501  29.255 38.627  31.13 38.627  31.13 36.752  33.004 36.752  33.004 34.878  34.879 34.878  34.879 33.003  36.753 33.003  36.753 31.129  38.628 31.129  38.628 29.254  40.502 29.254  40.502 27.38  42.377 27.38  42.377 25.505  44.251 25.505  44.251 23.631  46.126 23.631  46.126 21.756  48 21.756 ;
  END
END RIIO_BUMP_SNAG180_GND

MACRO RIIO_BUMP_SNAG180_PWR
  CLASS COVER ;
  ORIGIN 48 48 ;
  FOREIGN RIIO_BUMP_SNAG180_PWR -48 -48 ;
  SIZE 96 BY 96 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 1.026 -21.441 48 21.441 ;
        RECT 1.026 -25.5 44.882 25.5 ;
        RECT 1.026 -30.5 39.882 30.5 ;
        RECT 1.026 -35.5 34.882 35.5 ;
        RECT 1.026 -40.5 29.882 40.5 ;
        RECT 1.026 -45.5 24.882 45.5 ;
        RECT -19.882 -8.974 19.882 48 ;
        RECT -19.882 -48 19.882 -11.026 ;
        RECT -48 -22.382 -1.026 22.382 ;
        RECT -23 -46.441 -1.026 46.441 ;
        RECT -28 -42.382 -1.026 42.382 ;
        RECT -33 -37.382 -1.026 37.382 ;
        RECT -38 -32.382 -1.026 32.382 ;
        RECT -43 -27.382 -1.026 27.382 ;
    END
  END VDD
  OBS
    LAYER LB ;
      RECT -19.882 -48 19.882 48 ;
      RECT -21.441 -47.221 19.882 47.221 ;
      RECT -21.441 -46.75 22.382 46.75 ;
      RECT -23 -46.441 22.382 46.441 ;
      RECT -23 -45.5 24.882 45.5 ;
      RECT -25.5 -43.632 24.882 43.632 ;
      RECT -28 -42.382 24.882 42.382 ;
      RECT -28 -41.75 27.382 41.75 ;
      RECT -28 -40.5 29.882 40.5 ;
      RECT -30.5 -38.632 29.882 38.632 ;
      RECT -33 -37.382 29.882 37.382 ;
      RECT -33 -36.75 32.382 36.75 ;
      RECT -33 -35.5 34.882 35.5 ;
      RECT -35.5 -33.632 34.882 33.632 ;
      RECT -38 -32.382 34.882 32.382 ;
      RECT -38 -31.75 37.382 31.75 ;
      RECT -38 -30.5 39.882 30.5 ;
      RECT -40.5 -28.632 39.882 28.632 ;
      RECT -43 -27.382 39.882 27.382 ;
      RECT -43 -26.75 42.382 26.75 ;
      RECT -43 -25.5 44.882 25.5 ;
      RECT -45.5 -23.632 44.882 23.632 ;
      RECT -48 -22.382 44.882 22.382 ;
      RECT -48 -22.221 46.441 22.221 ;
      RECT -48 -21.441 48 21.441 ;
    LAYER VV ;
      RECT -19.261 -46.5 19.261 46.5 ;
      RECT -21.5 -45.381 19.261 45.381 ;
      RECT -21.5 -44 24.261 44 ;
      RECT -26.5 -41.761 24.261 41.761 ;
      RECT -26.5 -39 29.261 39 ;
      RECT -31.5 -36.761 29.261 36.761 ;
      RECT -31.5 -34 34.261 34 ;
      RECT -36.5 -31.761 34.261 31.761 ;
      RECT -36.5 -29 39.261 29 ;
      RECT -41.5 -26.761 39.261 26.761 ;
      RECT -41.5 -24 44.261 24 ;
      RECT -46.5 -21.761 44.261 21.761 ;
      RECT -46.5 -20.381 46.5 20.381 ;
    LAYER OVERLAP ;
      POLYGON  48 -21.757  46.125 -21.757  46.125 -23.632  44.25 -23.632  44.25 -25.506  42.376 -25.506  42.376 -27.381  40.501 -27.381  40.501 -29.255  38.627 -29.255  38.627 -31.13  36.752 -31.13  36.752 -33.004  34.878 -33.004  34.878 -34.879  33.003 -34.879  33.003 -36.753  31.129 -36.753  31.129 -38.628  29.254 -38.628  29.254 -40.502  27.38 -40.502  27.38 -42.377  25.505 -42.377  25.505 -44.251  23.631 -44.251  23.631 -46.126  21.756 -46.126  21.756 -48  -21.757 -48  -21.757 -46.125  -23.632 -46.125  -23.632 -44.25  -25.506 -44.25  -25.506 -42.376  -27.381 -42.376  -27.381 -40.501  -29.255 -40.501  -29.255 -38.627  -31.13 -38.627  -31.13 -36.752  -33.004 -36.752  -33.004 -34.878  -34.879 -34.878  -34.879 -33.003  -36.753 -33.003  -36.753 -31.129  -38.628 -31.129  -38.628 -29.254  -40.502 -29.254  -40.502 -27.38  -42.377 -27.38  -42.377 -25.505  -44.251 -25.505  -44.251 -23.631  -46.126 -23.631  -46.126 -21.756  -48 -21.756  -48 21.757  -46.125 21.757  -46.125 23.632  -44.25 23.632  -44.25 25.506  -42.376 25.506  -42.376 27.381  -40.501 27.381  -40.501 29.255  -38.627 29.255  -38.627 31.13  -36.752 31.13  -36.752 33.004  -34.878 33.004  -34.878 34.879  -33.003 34.879  -33.003 36.753  -31.129 36.753  -31.129 38.628  -29.254 38.628  -29.254 40.502  -27.38 40.502  -27.38 42.377  -25.505 42.377  -25.505 44.251  -23.631 44.251  -23.631 46.126  -21.756 46.126  -21.756 48  21.757 48  21.757 46.125  23.632 46.125  23.632 44.25  25.506 44.25  25.506 42.376  27.381 42.376  27.381 40.501  29.255 40.501  29.255 38.627  31.13 38.627  31.13 36.752  33.004 36.752  33.004 34.878  34.879 34.878  34.879 33.003  36.753 33.003  36.753 31.129  38.628 31.129  38.628 29.254  40.502 29.254  40.502 27.38  42.377 27.38  42.377 25.505  44.251 25.505  44.251 23.631  46.126 23.631  46.126 21.756  48 21.756 ;
  END
END RIIO_BUMP_SNAG180_PWR

MACRO RIIO_BUMP_SNAG180_SIG
  CLASS COVER ;
  ORIGIN 48 48 ;
  FOREIGN RIIO_BUMP_SNAG180_SIG -48 -48 ;
  SIZE 96 BY 96 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.210704 LAYER LB ;
    PORT
      LAYER LB ;
        RECT 1.026 -21.441 48 21.441 ;
        RECT 1.026 -25.5 44.882 25.5 ;
        RECT 1.026 -30.5 39.882 30.5 ;
        RECT 1.026 -35.5 34.882 35.5 ;
        RECT 1.026 -40.5 29.882 40.5 ;
        RECT 1.026 -45.5 24.882 45.5 ;
        RECT -19.882 -8.974 19.882 48 ;
        RECT -19.882 -48 19.882 -11.026 ;
        RECT -48 -22.382 -1.026 22.382 ;
        RECT -23 -46.441 -1.026 46.441 ;
        RECT -28 -42.382 -1.026 42.382 ;
        RECT -33 -37.382 -1.026 37.382 ;
        RECT -38 -32.382 -1.026 32.382 ;
        RECT -43 -27.382 -1.026 27.382 ;
    END
  END PAD
  OBS
    LAYER LB ;
      RECT -19.882 -48 19.882 48 ;
      RECT -21.441 -47.221 19.882 47.221 ;
      RECT -21.441 -46.75 22.382 46.75 ;
      RECT -23 -46.441 22.382 46.441 ;
      RECT -23 -45.5 24.882 45.5 ;
      RECT -25.5 -43.632 24.882 43.632 ;
      RECT -28 -42.382 24.882 42.382 ;
      RECT -28 -41.75 27.382 41.75 ;
      RECT -28 -40.5 29.882 40.5 ;
      RECT -30.5 -38.632 29.882 38.632 ;
      RECT -33 -37.382 29.882 37.382 ;
      RECT -33 -36.75 32.382 36.75 ;
      RECT -33 -35.5 34.882 35.5 ;
      RECT -35.5 -33.632 34.882 33.632 ;
      RECT -38 -32.382 34.882 32.382 ;
      RECT -38 -31.75 37.382 31.75 ;
      RECT -38 -30.5 39.882 30.5 ;
      RECT -40.5 -28.632 39.882 28.632 ;
      RECT -43 -27.382 39.882 27.382 ;
      RECT -43 -26.75 42.382 26.75 ;
      RECT -43 -25.5 44.882 25.5 ;
      RECT -45.5 -23.632 44.882 23.632 ;
      RECT -48 -22.382 44.882 22.382 ;
      RECT -48 -22.221 46.441 22.221 ;
      RECT -48 -21.441 48 21.441 ;
    LAYER VV ;
      RECT -19.261 -46.5 19.261 46.5 ;
      RECT -21.5 -45.381 19.261 45.381 ;
      RECT -21.5 -44 24.261 44 ;
      RECT -26.5 -41.761 24.261 41.761 ;
      RECT -26.5 -39 29.261 39 ;
      RECT -31.5 -36.761 29.261 36.761 ;
      RECT -31.5 -34 34.261 34 ;
      RECT -36.5 -31.761 34.261 31.761 ;
      RECT -36.5 -29 39.261 29 ;
      RECT -41.5 -26.761 39.261 26.761 ;
      RECT -41.5 -24 44.261 24 ;
      RECT -46.5 -21.761 44.261 21.761 ;
      RECT -46.5 -20.381 46.5 20.381 ;
    LAYER OVERLAP ;
      POLYGON  48 -21.757  46.125 -21.757  46.125 -23.632  44.25 -23.632  44.25 -25.506  42.376 -25.506  42.376 -27.381  40.501 -27.381  40.501 -29.255  38.627 -29.255  38.627 -31.13  36.752 -31.13  36.752 -33.004  34.878 -33.004  34.878 -34.879  33.003 -34.879  33.003 -36.753  31.129 -36.753  31.129 -38.628  29.254 -38.628  29.254 -40.502  27.38 -40.502  27.38 -42.377  25.505 -42.377  25.505 -44.251  23.631 -44.251  23.631 -46.126  21.756 -46.126  21.756 -48  -21.757 -48  -21.757 -46.125  -23.632 -46.125  -23.632 -44.25  -25.506 -44.25  -25.506 -42.376  -27.381 -42.376  -27.381 -40.501  -29.255 -40.501  -29.255 -38.627  -31.13 -38.627  -31.13 -36.752  -33.004 -36.752  -33.004 -34.878  -34.879 -34.878  -34.879 -33.003  -36.753 -33.003  -36.753 -31.129  -38.628 -31.129  -38.628 -29.254  -40.502 -29.254  -40.502 -27.38  -42.377 -27.38  -42.377 -25.505  -44.251 -25.505  -44.251 -23.631  -46.126 -23.631  -46.126 -21.756  -48 -21.756  -48 21.757  -46.125 21.757  -46.125 23.632  -44.25 23.632  -44.25 25.506  -42.376 25.506  -42.376 27.381  -40.501 27.381  -40.501 29.255  -38.627 29.255  -38.627 31.13  -36.752 31.13  -36.752 33.004  -34.878 33.004  -34.878 34.879  -33.003 34.879  -33.003 36.753  -31.129 36.753  -31.129 38.628  -29.254 38.628  -29.254 40.502  -27.38 40.502  -27.38 42.377  -25.505 42.377  -25.505 44.251  -23.631 44.251  -23.631 46.126  -21.756 46.126  -21.756 48  21.757 48  21.757 46.125  23.632 46.125  23.632 44.25  25.506 44.25  25.506 42.376  27.381 42.376  27.381 40.501  29.255 40.501  29.255 38.627  31.13 38.627  31.13 36.752  33.004 36.752  33.004 34.878  34.879 34.878  34.879 33.003  36.753 33.003  36.753 31.129  38.628 31.129  38.628 29.254  40.502 29.254  40.502 27.38  42.377 27.38  42.377 25.505  44.251 25.505  44.251 23.631  46.126 23.631  46.126 21.756  48 21.756 ;
  END
END RIIO_BUMP_SNAG180_SIG

MACRO RIIO_BOND20x10_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND20x10_INNER_GND 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 10.01 0 29.99 10 ;
      LAYER QB ;
        RECT 15 0 25 10 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 10 5 29.99 10 ;
      RECT 10.01 0 30 5 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER JV ;
      RECT 0 0 40 10 ;
    LAYER YS ;
      RECT 0 0 40 10 ;
    LAYER JW ;
      RECT 0 0 40 10 ;
    LAYER QB ;
      RECT 0 0 40 10 ;
    LAYER QA ;
      RECT 0 0 40 10 ;
    LAYER JA ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND20x10_INNER_GND

MACRO RIIO_BOND20x10_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND20x10_INNER_PWR 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 10 0 30 10 ;
      LAYER QB ;
        RECT 15 0 25 10 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 10 0 30 10 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER JV ;
      RECT 0 0 40 10 ;
    LAYER YS ;
      RECT 0 0 40 10 ;
    LAYER JW ;
      RECT 0 0 40 10 ;
    LAYER QB ;
      RECT 0 0 40 10 ;
    LAYER QA ;
      RECT 0 0 40 10 ;
    LAYER JA ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND20x10_INNER_PWR

MACRO RIIO_BOND20x10_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND20x10_INNER_SIG 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 175 LAYER QB ;
    ANTENNAPARTIALCUTAREA 43.74 LAYER VV ;
    PORT
      LAYER QB ;
        RECT 15 0 25 10 ;
      LAYER LB ;
        RECT 10 0 30 10 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 10 0 30 10 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER JV ;
      RECT 0 0 40 10 ;
    LAYER YS ;
      RECT 0 0 40 10 ;
    LAYER JW ;
      RECT 0 0 40 10 ;
    LAYER QB ;
      RECT 0 0 40 10 ;
    LAYER QA ;
      RECT 0 0 40 10 ;
    LAYER JA ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND20x10_INNER_SIG

MACRO RIIO_BOND60_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_INNER_GND 0 0 ;
  SIZE 60 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 10 0 50 70 ;
      LAYER QB ;
        RECT 10 69 50 70 ;
      LAYER QA ;
        RECT 10 69 50 70 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER JV ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER YS ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER JW ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER QB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER QA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER JA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  50 60  50 70  10 70  10 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_INNER_GND

MACRO RIIO_BOND60_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_INNER_PWR 0 0 ;
  SIZE 60 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 10 0 50 70 ;
      LAYER QB ;
        RECT 10 69 50 70 ;
      LAYER QA ;
        RECT 10 69 50 70 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER JV ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER YS ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER JW ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER QB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER QA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER JA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  50 60  50 70  10 70  10 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_INNER_PWR

MACRO RIIO_BOND60_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_INNER_SIG 0 0 ;
  SIZE 60 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2635 LAYER QA ;
    ANTENNAPARTIALMETALAREA 2809.16 LAYER QB ;
    ANTENNAPARTIALCUTAREA 616.32 LAYER JW ;
    ANTENNAPARTIALCUTAREA 422.82 LAYER VV ;
    PORT
      LAYER QA ;
        RECT 10 69 50 70 ;
      LAYER QB ;
        RECT 10 69 50 70 ;
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 10 0 50 70 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER JV ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER YS ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER JW ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER QB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER QA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER JA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  50 60  50 70  10 70  10 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_INNER_SIG

MACRO RIIO_BOND60_OUTER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_OUTER_GND 0 0 ;
  SIZE 60 BY 140 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 12.5 0 47.5 140 ;
      LAYER QB ;
        RECT 12.5 139 47.5 140 ;
      LAYER QA ;
        RECT 12.5 139 47.5 140 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER JV ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER YS ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER JW ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER QB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER QA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER JA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  47.5 60  47.5 140  12.5 140  12.5 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_OUTER_GND

MACRO RIIO_BOND60_OUTER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_OUTER_PWR 0 0 ;
  SIZE 60 BY 140 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 12.5 0 47.5 140 ;
      LAYER QB ;
        RECT 12.5 139 47.5 140 ;
      LAYER QA ;
        RECT 12.5 139 47.5 140 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER JV ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER YS ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER JW ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER QB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER QA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER JA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  47.5 60  47.5 140  12.5 140  12.5 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_OUTER_PWR

MACRO RIIO_BOND60_OUTER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_OUTER_SIG 0 0 ;
  SIZE 60 BY 140 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4540 LAYER QA ;
    ANTENNAPARTIALMETALAREA 4689.16 LAYER QB ;
    ANTENNAPARTIALCUTAREA 1054.08 LAYER JW ;
    ANTENNAPARTIALCUTAREA 816.48 LAYER VV ;
    PORT
      LAYER QA ;
        RECT 12.5 139 47.5 140 ;
      LAYER QB ;
        RECT 12.5 139 47.5 140 ;
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 12.5 0 47.5 140 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER JV ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER YS ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER JW ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER QB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER QA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER JA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  47.5 60  47.5 140  12.5 140  12.5 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_OUTER_SIG

MACRO RIIO_BOND60_PLAIN_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_PLAIN_GND 0 0 ;
  SIZE 60 BY 60 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 0 0 60 60 ;
    LAYER JV ;
      RECT 0 0 60 60 ;
    LAYER YS ;
      RECT 0 0 60 60 ;
    LAYER JW ;
      RECT 0 0 60 60 ;
    LAYER QB ;
      RECT 0 0 60 60 ;
    LAYER QA ;
      RECT 0 0 60 60 ;
    LAYER JA ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 0 0 60 60 ;
  END
END RIIO_BOND60_PLAIN_GND

MACRO RIIO_BOND60_PLAIN_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_PLAIN_PWR 0 0 ;
  SIZE 60 BY 60 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 0 0 60 60 ;
    LAYER JV ;
      RECT 0 0 60 60 ;
    LAYER YS ;
      RECT 0 0 60 60 ;
    LAYER JW ;
      RECT 0 0 60 60 ;
    LAYER QB ;
      RECT 0 0 60 60 ;
    LAYER QA ;
      RECT 0 0 60 60 ;
    LAYER JA ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 0 0 60 60 ;
  END
END RIIO_BOND60_PLAIN_PWR

MACRO RIIO_BOND60_PLAIN_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_PLAIN_SIG 0 0 ;
  SIZE 60 BY 60 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 0 0 60 60 ;
    LAYER JV ;
      RECT 0 0 60 60 ;
    LAYER YS ;
      RECT 0 0 60 60 ;
    LAYER JW ;
      RECT 0 0 60 60 ;
    LAYER QB ;
      RECT 0 0 60 60 ;
    LAYER QA ;
      RECT 0 0 60 60 ;
    LAYER JA ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 0 0 60 60 ;
  END
END RIIO_BOND60_PLAIN_SIG

MACRO RIIO_BOND60x90_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_GND 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
      LAYER QB ;
        RECT 10 99 50 100 ;
      LAYER QA ;
        RECT 10 99 50 100 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_GND

MACRO RIIO_BOND60x90_INNER_GND_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_GND_CESD 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
      LAYER QB ;
        RECT 10 99 50 100 ;
      LAYER QA ;
        RECT 10 99 50 100 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_GND_CESD

MACRO RIIO_BOND60x90_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_PWR 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
      LAYER QB ;
        RECT 10 99 50 100 ;
      LAYER QA ;
        RECT 10 99 50 100 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_PWR

MACRO RIIO_BOND60x90_INNER_PWR_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_PWR_CESD 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
      LAYER QB ;
        RECT 10 99 50 100 ;
      LAYER QA ;
        RECT 10 99 50 100 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_PWR_CESD

MACRO RIIO_BOND60x90_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_SIG 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3910 LAYER QA ;
    ANTENNAPARTIALMETALAREA 4117.16 LAYER QB ;
    ANTENNAPARTIALCUTAREA 910.08 LAYER JW ;
    ANTENNAPARTIALCUTAREA 510.3 LAYER VV ;
    PORT
      LAYER QA ;
        RECT 10 99 50 100 ;
      LAYER QB ;
        RECT 10 99 50 100 ;
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_SIG

MACRO RIIO_BOND60x90_INNER_SIG_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_SIG_CESD 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3910 LAYER QA ;
    ANTENNAPARTIALMETALAREA 4117.16 LAYER QB ;
    ANTENNAPARTIALCUTAREA 910.08 LAYER JW ;
    ANTENNAPARTIALCUTAREA 510.3 LAYER VV ;
    PORT
      LAYER QA ;
        RECT 10 99 50 100 ;
      LAYER QB ;
        RECT 10 99 50 100 ;
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_SIG_CESD

MACRO RIIO_BOND60x90_OUTER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_GND 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
      LAYER QB ;
        RECT 12.5 199 47.5 200 ;
      LAYER QA ;
        RECT 12.5 199 47.5 200 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_GND

MACRO RIIO_BOND60x90_OUTER_GND_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_GND_CESD 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
      LAYER QB ;
        RECT 12.5 199 47.5 200 ;
      LAYER QA ;
        RECT 12.5 199 47.5 200 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_GND_CESD

MACRO RIIO_BOND60x90_OUTER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_PWR 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
      LAYER QB ;
        RECT 12.5 199 47.5 200 ;
      LAYER QA ;
        RECT 12.5 199 47.5 200 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_PWR

MACRO RIIO_BOND60x90_OUTER_PWR_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_PWR_CESD 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
      LAYER QB ;
        RECT 12.5 199 47.5 200 ;
      LAYER QA ;
        RECT 12.5 199 47.5 200 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_PWR_CESD

MACRO RIIO_BOND60x90_OUTER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_SIG 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6640 LAYER QA ;
    ANTENNAPARTIALMETALAREA 6822.16 LAYER QB ;
    ANTENNAPARTIALCUTAREA 1537.92 LAYER JW ;
    ANTENNAPARTIALCUTAREA 1078.92 LAYER VV ;
    PORT
      LAYER QA ;
        RECT 12.5 199 47.5 200 ;
      LAYER QB ;
        RECT 12.5 199 47.5 200 ;
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_SIG

MACRO RIIO_BOND60x90_OUTER_SIG_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_SIG_CESD 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6640 LAYER QA ;
    ANTENNAPARTIALMETALAREA 6822.16 LAYER QB ;
    ANTENNAPARTIALCUTAREA 1537.92 LAYER JW ;
    ANTENNAPARTIALCUTAREA 1078.92 LAYER VV ;
    PORT
      LAYER QA ;
        RECT 12.5 199 47.5 200 ;
      LAYER QB ;
        RECT 12.5 199 47.5 200 ;
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_SIG_CESD

MACRO RIIO_BOND60x90_PLAIN_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_GND 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_GND

MACRO RIIO_BOND60x90_PLAIN_GND_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_GND_CESD 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_GND_CESD

MACRO RIIO_BOND60x90_PLAIN_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_PWR 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_PWR

MACRO RIIO_BOND60x90_PLAIN_PWR_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_PWR_CESD 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_PWR_CESD

MACRO RIIO_BOND60x90_PLAIN_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_SIG 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_SIG

MACRO RIIO_BOND60x90_PLAIN_SIG_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_SIG_CESD 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER JV ;
      RECT 0 0 60 90 ;
    LAYER YS ;
      RECT 0 0 60 90 ;
    LAYER JW ;
      RECT 0 0 60 90 ;
    LAYER QB ;
      RECT 0 0 60 90 ;
    LAYER QA ;
      RECT 0 0 60 90 ;
    LAYER JA ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_SIG_CESD

MACRO RIIO_BOND64_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_INNER_GND 0 0 ;
  SIZE 64 BY 72 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 12 0 52 72 ;
      LAYER QB ;
        RECT 12 71 52 72 ;
      LAYER QA ;
        RECT 12 71 52 72 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER JV ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER YS ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER JW ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER QB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER QA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER JA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 72  12 72  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_INNER_GND

MACRO RIIO_BOND64_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_INNER_PWR 0 0 ;
  SIZE 64 BY 72 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 12 0 52 72 ;
      LAYER QB ;
        RECT 12 71 52 72 ;
      LAYER QA ;
        RECT 12 71 52 72 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER JV ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER YS ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER JW ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER QB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER QA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER JA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 72  12 72  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_INNER_PWR

MACRO RIIO_BOND64_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_INNER_SIG 0 0 ;
  SIZE 64 BY 72 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2529.6 LAYER QA ;
    ANTENNAPARTIALMETALAREA 2807.84 LAYER QB ;
    ANTENNAPARTIALCUTAREA 270.72 LAYER JW ;
    ANTENNAPARTIALCUTAREA 408.24 LAYER VV ;
    PORT
      LAYER QA ;
        RECT 12 71 52 72 ;
      LAYER QB ;
        RECT 12 71 52 72 ;
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 12 0 52 72 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER JV ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER YS ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER JW ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER QB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER QA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER JA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 72  12 72  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_INNER_SIG

MACRO RIIO_BOND64_OUTER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_OUTER_GND 0 0 ;
  SIZE 64 BY 144 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 11.998 0 52 144 ;
      LAYER QB ;
        RECT 12 143 52 144 ;
      LAYER QA ;
        RECT 12 143 52 144 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 11.998 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER JV ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER YS ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER JW ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER QB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER QA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER JA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 144  12 144  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_OUTER_GND

MACRO RIIO_BOND64_OUTER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_OUTER_PWR 0 0 ;
  SIZE 64 BY 144 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 11.998 0 52 144 ;
      LAYER QB ;
        RECT 12 143 52 144 ;
      LAYER QA ;
        RECT 12 143 52 144 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 11.998 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER JV ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER YS ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER JW ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER QB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER QA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER JA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 144  12 144  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_OUTER_PWR

MACRO RIIO_BOND64_OUTER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_OUTER_SIG 0 0 ;
  SIZE 64 BY 144 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4152 LAYER QA ;
    ANTENNAPARTIALMETALAREA 4190.24 LAYER QB ;
    ANTENNAPARTIALCUTAREA 466.56 LAYER JW ;
    ANTENNAPARTIALCUTAREA 816.48 LAYER VV ;
    PORT
      LAYER QA ;
        RECT 12 143 52 144 ;
      LAYER QB ;
        RECT 12 143 52 144 ;
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 11.998 0 52 144 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 11.998 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER JV ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER YS ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER JW ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER QB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER QA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER JA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 144  12 144  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_OUTER_SIG

MACRO RIIO_BOND64_PLAIN_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_PLAIN_GND 0 0 ;
  SIZE 64 BY 64 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 0 0 64 64 ;
    LAYER JV ;
      RECT 0 0 64 64 ;
    LAYER YS ;
      RECT 0 0 64 64 ;
    LAYER JW ;
      RECT 0 0 64 64 ;
    LAYER QB ;
      RECT 0 0 64 64 ;
    LAYER QA ;
      RECT 0 0 64 64 ;
    LAYER JA ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 0 0 64 64 ;
  END
END RIIO_BOND64_PLAIN_GND

MACRO RIIO_BOND64_PLAIN_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_PLAIN_PWR 0 0 ;
  SIZE 64 BY 64 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 0 0 64 64 ;
    LAYER JV ;
      RECT 0 0 64 64 ;
    LAYER YS ;
      RECT 0 0 64 64 ;
    LAYER JW ;
      RECT 0 0 64 64 ;
    LAYER QB ;
      RECT 0 0 64 64 ;
    LAYER QA ;
      RECT 0 0 64 64 ;
    LAYER JA ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 0 0 64 64 ;
  END
END RIIO_BOND64_PLAIN_PWR

MACRO RIIO_BOND64_PLAIN_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_PLAIN_SIG 0 0 ;
  SIZE 64 BY 64 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 0 0 64 64 ;
    LAYER JV ;
      RECT 0 0 64 64 ;
    LAYER YS ;
      RECT 0 0 64 64 ;
    LAYER JW ;
      RECT 0 0 64 64 ;
    LAYER QB ;
      RECT 0 0 64 64 ;
    LAYER QA ;
      RECT 0 0 64 64 ;
    LAYER JA ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 0 0 64 64 ;
  END
END RIIO_BOND64_PLAIN_SIG

MACRO RIIO_BOND70_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_INNER_GND 0 0 ;
  SIZE 70 BY 80 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 15 0 55 80 ;
      LAYER QB ;
        RECT 15 79 55 80 ;
      LAYER QA ;
        RECT 15 79 55 80 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER JV ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER YS ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER JW ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER QB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER QA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER JA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  55 70  55 80  15 80  15 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_INNER_GND

MACRO RIIO_BOND70_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_INNER_PWR 0 0 ;
  SIZE 70 BY 80 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 15 0 55 80 ;
      LAYER QB ;
        RECT 15 79 55 80 ;
      LAYER QA ;
        RECT 15 79 55 80 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER JV ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER YS ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER JW ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER QB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER QA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER JA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  55 70  55 80  15 80  15 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_INNER_PWR

MACRO RIIO_BOND70_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_INNER_SIG 0 0 ;
  SIZE 70 BY 80 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3560 LAYER QA ;
    ANTENNAPARTIALMETALAREA 3585 LAYER QB ;
    ANTENNAPARTIALCUTAREA 829.44 LAYER JW ;
    ANTENNAPARTIALCUTAREA 481.14 LAYER VV ;
    PORT
      LAYER QA ;
        RECT 15 79 55 80 ;
      LAYER QB ;
        RECT 15 79 55 80 ;
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 15 0 55 80 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER JV ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER YS ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER JW ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER QB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER QA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER JA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  55 70  55 80  15 80  15 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_INNER_SIG

MACRO RIIO_BOND70_OUTER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_OUTER_GND 0 0 ;
  SIZE 70 BY 160 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 17.5 0 52.5 160 ;
      LAYER QB ;
        RECT 17.5 159 52.5 160 ;
      LAYER QA ;
        RECT 17.5 159 52.5 160 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER JV ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER YS ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER JW ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER QB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER QA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER JA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  52.5 70  52.5 160  17.5 160  17.5 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_OUTER_GND

MACRO RIIO_BOND70_OUTER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_OUTER_PWR 0 0 ;
  SIZE 70 BY 160 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 17.5 0 52.5 160 ;
      LAYER QB ;
        RECT 17.5 159 52.5 160 ;
      LAYER QA ;
        RECT 17.5 159 52.5 160 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER JV ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER YS ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER JW ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER QB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER QA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER JA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  52.5 70  52.5 160  17.5 160  17.5 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_OUTER_PWR

MACRO RIIO_BOND70_OUTER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_OUTER_SIG 0 0 ;
  SIZE 70 BY 160 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5740 LAYER QA ;
    ANTENNAPARTIALMETALAREA 5740 LAYER QB ;
    ANTENNAPARTIALCUTAREA 1330.56 LAYER JW ;
    ANTENNAPARTIALCUTAREA 933.12 LAYER VV ;
    PORT
      LAYER QA ;
        RECT 17.5 159 52.5 160 ;
      LAYER QB ;
        RECT 17.5 159 52.5 160 ;
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 17.5 0 52.5 160 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER JV ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER YS ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER JW ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER QB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER QA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER JA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  52.5 70  52.5 160  17.5 160  17.5 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_OUTER_SIG

MACRO RIIO_BOND70_PLAIN_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_PLAIN_GND 0 0 ;
  SIZE 70 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 0 0 70 70 ;
    LAYER JV ;
      RECT 0 0 70 70 ;
    LAYER YS ;
      RECT 0 0 70 70 ;
    LAYER JW ;
      RECT 0 0 70 70 ;
    LAYER QB ;
      RECT 0 0 70 70 ;
    LAYER QA ;
      RECT 0 0 70 70 ;
    LAYER JA ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 0 0 70 70 ;
  END
END RIIO_BOND70_PLAIN_GND

MACRO RIIO_BOND70_PLAIN_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_PLAIN_PWR 0 0 ;
  SIZE 70 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 0 0 70 70 ;
    LAYER JV ;
      RECT 0 0 70 70 ;
    LAYER YS ;
      RECT 0 0 70 70 ;
    LAYER JW ;
      RECT 0 0 70 70 ;
    LAYER QB ;
      RECT 0 0 70 70 ;
    LAYER QA ;
      RECT 0 0 70 70 ;
    LAYER JA ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 0 0 70 70 ;
  END
END RIIO_BOND70_PLAIN_PWR

MACRO RIIO_BOND70_PLAIN_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_PLAIN_SIG 0 0 ;
  SIZE 70 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 0 0 70 70 ;
    LAYER JV ;
      RECT 0 0 70 70 ;
    LAYER YS ;
      RECT 0 0 70 70 ;
    LAYER JW ;
      RECT 0 0 70 70 ;
    LAYER QB ;
      RECT 0 0 70 70 ;
    LAYER QA ;
      RECT 0 0 70 70 ;
    LAYER JA ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 0 0 70 70 ;
  END
END RIIO_BOND70_PLAIN_SIG

MACRO RIIO_BOND80x100_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_INNER_GND 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT -20 -110 60 -10 ;
        RECT 0 -110 40 10 ;
      LAYER QB ;
        RECT 15 0 25 10 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 0 -110 40 10 ;
      RECT -20 -110 60 -10 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER JV ;
      RECT 0 0 40 10 ;
    LAYER YS ;
      RECT 0 0 40 10 ;
    LAYER JW ;
      RECT 0 0 40 10 ;
    LAYER QB ;
      RECT 0 0 40 10 ;
    LAYER QA ;
      RECT 0 0 40 10 ;
    LAYER JA ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND80x100_INNER_GND

MACRO RIIO_BOND80x100_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_INNER_PWR 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT -20 -110 60 -10 ;
        RECT 0 -110 40 10 ;
      LAYER QB ;
        RECT 15 0 25 10 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 0 -110 40 10 ;
      RECT -20 -110 60 -10 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER JV ;
      RECT 0 0 40 10 ;
    LAYER YS ;
      RECT 0 0 40 10 ;
    LAYER JW ;
      RECT 0 0 40 10 ;
    LAYER QB ;
      RECT 0 0 40 10 ;
    LAYER QA ;
      RECT 0 0 40 10 ;
    LAYER JA ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND80x100_INNER_PWR

MACRO RIIO_BOND80x100_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_INNER_SIG 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 225 LAYER QB ;
    ANTENNAPARTIALCUTAREA 72.9 LAYER VV ;
    PORT
      LAYER QB ;
        RECT 15 0 25 10 ;
      LAYER LB ;
        RECT -20 -110 60 -10 ;
        RECT 0 -110 40 10 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 0 -110 40 10 ;
      RECT -20 -110 60 -10 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER JV ;
      RECT 0 0 40 10 ;
    LAYER YS ;
      RECT 0 0 40 10 ;
    LAYER JW ;
      RECT 0 0 40 10 ;
    LAYER QB ;
      RECT 0 0 40 10 ;
    LAYER QA ;
      RECT 0 0 40 10 ;
    LAYER JA ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND80x100_INNER_SIG

MACRO RIIO_BOND80x100_PLAIN_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_PLAIN_GND 0 0 ;
  SIZE 80 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 80 100 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 100 ;
    LAYER M1 ;
      RECT 0 0 80 100 ;
    LAYER V1 ;
      RECT 0 0 80 100 ;
    LAYER M2 ;
      RECT 0 0 80 100 ;
    LAYER A1 ;
      RECT 0 0 80 100 ;
    LAYER C2 ;
      RECT 0 0 80 100 ;
    LAYER LB ;
      RECT 0 0 80 100 ;
    LAYER VV ;
      RECT 0 0 80 100 ;
    LAYER CB ;
      RECT 0 0 80 100 ;
    LAYER JV ;
      RECT 0 0 80 100 ;
    LAYER YS ;
      RECT 0 0 80 100 ;
    LAYER JW ;
      RECT 0 0 80 100 ;
    LAYER QB ;
      RECT 0 0 80 100 ;
    LAYER QA ;
      RECT 0 0 80 100 ;
    LAYER JA ;
      RECT 0 0 80 100 ;
    LAYER AY ;
      RECT 0 0 80 100 ;
    LAYER C1 ;
      RECT 0 0 80 100 ;
    LAYER C5 ;
      RECT 0 0 80 100 ;
    LAYER C4 ;
      RECT 0 0 80 100 ;
    LAYER C3 ;
      RECT 0 0 80 100 ;
    LAYER A4 ;
      RECT 0 0 80 100 ;
    LAYER A3 ;
      RECT 0 0 80 100 ;
    LAYER A2 ;
      RECT 0 0 80 100 ;
  END
END RIIO_BOND80x100_PLAIN_GND

MACRO RIIO_BOND80x100_PLAIN_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_PLAIN_PWR 0 0 ;
  SIZE 80 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 80 100 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 100 ;
    LAYER M1 ;
      RECT 0 0 80 100 ;
    LAYER V1 ;
      RECT 0 0 80 100 ;
    LAYER M2 ;
      RECT 0 0 80 100 ;
    LAYER A1 ;
      RECT 0 0 80 100 ;
    LAYER C2 ;
      RECT 0 0 80 100 ;
    LAYER LB ;
      RECT 0 0 80 100 ;
    LAYER VV ;
      RECT 0 0 80 100 ;
    LAYER CB ;
      RECT 0 0 80 100 ;
    LAYER JV ;
      RECT 0 0 80 100 ;
    LAYER YS ;
      RECT 0 0 80 100 ;
    LAYER JW ;
      RECT 0 0 80 100 ;
    LAYER QB ;
      RECT 0 0 80 100 ;
    LAYER QA ;
      RECT 0 0 80 100 ;
    LAYER JA ;
      RECT 0 0 80 100 ;
    LAYER AY ;
      RECT 0 0 80 100 ;
    LAYER C1 ;
      RECT 0 0 80 100 ;
    LAYER C5 ;
      RECT 0 0 80 100 ;
    LAYER C4 ;
      RECT 0 0 80 100 ;
    LAYER C3 ;
      RECT 0 0 80 100 ;
    LAYER A4 ;
      RECT 0 0 80 100 ;
    LAYER A3 ;
      RECT 0 0 80 100 ;
    LAYER A2 ;
      RECT 0 0 80 100 ;
  END
END RIIO_BOND80x100_PLAIN_PWR

MACRO RIIO_BOND80x100_PLAIN_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_PLAIN_SIG 0 0 ;
  SIZE 80 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 80 100 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 80 100 ;
    LAYER M1 ;
      RECT 0 0 80 100 ;
    LAYER V1 ;
      RECT 0 0 80 100 ;
    LAYER M2 ;
      RECT 0 0 80 100 ;
    LAYER A1 ;
      RECT 0 0 80 100 ;
    LAYER C2 ;
      RECT 0 0 80 100 ;
    LAYER LB ;
      RECT 0 0 80 100 ;
    LAYER VV ;
      RECT 0 0 80 100 ;
    LAYER CB ;
      RECT 0 0 80 100 ;
    LAYER JV ;
      RECT 0 0 80 100 ;
    LAYER YS ;
      RECT 0 0 80 100 ;
    LAYER JW ;
      RECT 0 0 80 100 ;
    LAYER QB ;
      RECT 0 0 80 100 ;
    LAYER QA ;
      RECT 0 0 80 100 ;
    LAYER JA ;
      RECT 0 0 80 100 ;
    LAYER AY ;
      RECT 0 0 80 100 ;
    LAYER C1 ;
      RECT 0 0 80 100 ;
    LAYER C5 ;
      RECT 0 0 80 100 ;
    LAYER C4 ;
      RECT 0 0 80 100 ;
    LAYER C3 ;
      RECT 0 0 80 100 ;
    LAYER A4 ;
      RECT 0 0 80 100 ;
    LAYER A3 ;
      RECT 0 0 80 100 ;
    LAYER A2 ;
      RECT 0 0 80 100 ;
  END
END RIIO_BOND80x100_PLAIN_SIG

END LIBRARY
