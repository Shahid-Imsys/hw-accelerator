-- PEC Part of NoC simulation pkg
-- 
-- Design: Imsys AB
-- Implemented: Bengt Andersson
-- Revision 0


library ieee;
use ieee.std_logic_1164.all;

library work;
use work.defines.all;



entity PEC is 
port (
	
);
end entity PEC;



architecture PEC_rtl of PEC is
begin

end architecture PEC_rtl;