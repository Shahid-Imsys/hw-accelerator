VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RIIO_EG1D80V_BIAS_RVT28_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_BIAS_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 59.35 60 62.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 64.05 60 67.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
    END
  END VDD
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.352 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 0 39.575 60 40.825 ;
    END
  END VBIAS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER OI ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      LAYER OI ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      LAYER OI ;
        RECT 54.05 0 57.65 58.25 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 58.25 ;
        RECT 35.25 0 38.85 58.25 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 58.25 ;
        RECT 11.75 0 15.35 58.25 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 58.25 ;
      LAYER IA ;
        RECT 0 3.67 60 6.55 ;
        RECT 0 17.05 60 20.65 ;
        RECT 0 26.45 60 30.05 ;
        RECT 0 40.55 60 44.15 ;
        RECT 0 45.25 60 48.85 ;
        RECT 0 54.65 60 58.25 ;
    END
  END VSSIO
  PIN TRIM_CURV_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.87128 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03808 LAYER C1 ;
      ANTENNAMAXAREACAR 81.406755 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 45.65 79.84 45.81 80 ;
    END
  END TRIM_CURV_I[4]
  PIN TRIM_CURV_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.86008 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03808 LAYER C1 ;
      ANTENNAMAXAREACAR 80.343407 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 45.13 79.84 45.29 80 ;
    END
  END TRIM_CURV_I[3]
  PIN TRIM_CURV_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.05888 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04704 LAYER C1 ;
      ANTENNAMAXAREACAR 70.193878 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 44.61 79.84 44.77 80 ;
    END
  END TRIM_CURV_I[2]
  PIN TRIM_CURV_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.16948 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.07392 LAYER C1 ;
      ANTENNAMAXAREACAR 50.562432 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 44.09 79.84 44.25 80 ;
    END
  END TRIM_CURV_I[1]
  PIN TRIM_CURV_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.67248 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1456 LAYER C1 ;
      ANTENNAMAXAREACAR 27.374176 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 43.57 79.84 43.73 80 ;
    END
  END TRIM_CURV_I[0]
  PIN BG_VALID_N_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.08032 LAYER C1 ;
    ANTENNADIFFAREA 0.1045 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.099 LAYER C1 ;
      ANTENNAMAXAREACAR 10.462518 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 25.11 79.84 25.27 80 ;
    END
  END BG_VALID_N_O
  PIN EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4424 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 58.141304 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 13.67 79.84 13.83 80 ;
    END
  END EN_I
  PIN VTMP_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.97008 LAYER C1 ;
    ANTENNADIFFAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.4 LAYER C1 ;
      ANTENNAMAXAREACAR 2.244581 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 18.09 79.84 18.25 80 ;
    END
  END VTMP_O
  PIN VBG_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.97008 LAYER C1 ;
    ANTENNADIFFAREA 0.32 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.4 LAYER C1 ;
      ANTENNAMAXAREACAR 2.553479 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.45 79.84 14.61 80 ;
    END
  END VBG_O
  PIN IBIAS_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.87 79.84 6.03 80 ;
    END
  END IBIAS_O[15]
  PIN TRIM_BIAS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4424 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 58.054348 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 28.23 79.84 28.39 80 ;
    END
  END TRIM_BIAS_I[3]
  PIN TRIM_BIAS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4424 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 58.166149 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 24.59 79.84 24.75 80 ;
    END
  END TRIM_BIAS_I[2]
  PIN TRIM_BIAS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4424 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 58.029503 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 17.31 79.84 17.47 80 ;
    END
  END TRIM_BIAS_I[1]
  PIN TRIM_BIAS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4424 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 58.27795 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 20.95 79.84 21.11 80 ;
    END
  END TRIM_BIAS_I[0]
  PIN IBIAS_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.13 79.84 6.29 80 ;
    END
  END IBIAS_O[14]
  PIN IBIAS_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.39 79.84 6.55 80 ;
    END
  END IBIAS_O[13]
  PIN IBIAS_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.65 79.84 6.81 80 ;
    END
  END IBIAS_O[12]
  PIN IBIAS_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.91 79.84 7.07 80 ;
    END
  END IBIAS_O[11]
  PIN IBIAS_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 7.17 79.84 7.33 80 ;
    END
  END IBIAS_O[10]
  PIN IBIAS_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 7.43 79.84 7.59 80 ;
    END
  END IBIAS_O[9]
  PIN IBIAS_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 7.69 79.84 7.85 80 ;
    END
  END IBIAS_O[8]
  PIN IBIAS_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 8.47 79.84 8.63 80 ;
    END
  END IBIAS_O[7]
  PIN IBIAS_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 8.73 79.84 8.89 80 ;
    END
  END IBIAS_O[6]
  PIN IBIAS_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 9.51 79.84 9.67 80 ;
    END
  END IBIAS_O[5]
  PIN IBIAS_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 9.77 79.84 9.93 80 ;
    END
  END IBIAS_O[4]
  PIN IBIAS_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.55 79.84 10.71 80 ;
    END
  END IBIAS_O[3]
  PIN IBIAS_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.81 79.84 10.97 80 ;
    END
  END IBIAS_O[2]
  PIN IBIAS_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 11.07 79.84 11.23 80 ;
    END
  END IBIAS_O[1]
  PIN IBIAS_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96528 LAYER C1 ;
    ANTENNADIFFAREA 0.088 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 11.33 79.84 11.49 80 ;
    END
  END IBIAS_O[0]
  PIN BG_STARTUP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.09808 LAYER C1 ;
    ANTENNADIFFAREA 0.2528 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.474 LAYER C1 ;
      ANTENNAMAXAREACAR 6.261814 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 23.03 79.84 23.19 80 ;
    END
  END BG_STARTUP_I
  PIN TRIM_VBG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.12288 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03808 LAYER C1 ;
      ANTENNAMAXAREACAR 87.244667 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.93 79.84 40.09 80 ;
    END
  END TRIM_VBG_I[4]
  PIN TRIM_VBG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.06168 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03808 LAYER C1 ;
      ANTENNAMAXAREACAR 85.637524 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.41 79.84 39.57 80 ;
    END
  END TRIM_VBG_I[3]
  PIN TRIM_VBG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.35008 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04704 LAYER C1 ;
      ANTENNAMAXAREACAR 76.697598 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.89 79.84 39.05 80 ;
    END
  END TRIM_VBG_I[2]
  PIN TRIM_VBG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.49428 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.07392 LAYER C1 ;
      ANTENNAMAXAREACAR 54.639236 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 38.37 79.84 38.53 80 ;
    END
  END TRIM_VBG_I[1]
  PIN TRIM_VBG_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7464 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1456 LAYER C1 ;
      ANTENNAMAXAREACAR 29.124725 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.85 79.84 38.01 80 ;
    END
  END TRIM_VBG_I[0]
  PIN EN_VBIAS_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4424 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 58.253106 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 10.03 79.84 10.19 80 ;
    END
  END EN_VBIAS_I
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER YZ ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER WT ;
      RECT 0 0 60 80 ;
    LAYER BA ;
      RECT 0 0 60 80 ;
    LAYER WA ;
      RECT 0 0 60 80 ;
    LAYER BB ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_BIAS_RVT28_V

MACRO RIIO_EG1D80V_GPIO_RVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPIO_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52912 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.704969 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.24 79.84 19.4 80 ;
    END
  END CO_I
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 400.1975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 135.895 LAYER BB ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER IA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 241.9675 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 15.4548 LAYER WA ;
    ANTENNAPARTIALCUTAREA 10.4976 LAYER WT ;
    ANTENNAPARTIALCUTAREA 13.226976 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A2 ;
    ANTENNADIFFAREA 208.5584 LAYER BA ;
    ANTENNADIFFAREA 208.5584 LAYER C3 ;
    ANTENNADIFFAREA 208.5584 LAYER BB ;
    ANTENNADIFFAREA 208.5584 LAYER IA ;
    ANTENNADIFFAREA 208.5584 LAYER OI ;
    ANTENNADIFFAREA 208.5584 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN DI_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.02096 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.78 79.84 39.94 80 ;
    END
  END DI_O[0]
  PIN DI_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.01968 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.96 79.84 38.12 80 ;
    END
  END DI_O[1]
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.76592 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.287798 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 8.32 79.84 8.48 80 ;
    END
  END DO_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7984 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.962733 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 24.18 79.84 24.34 80 ;
    END
  END DS_I[0]
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.796 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.829193 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 26.78 79.84 26.94 80 ;
    END
  END DS_I[1]
  PIN DS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53232 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 140.512422 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 9.62 79.84 9.78 80 ;
    END
  END DS_I[2]
  PIN DS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52864 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.773292 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 3.9 79.84 4.06 80 ;
    END
  END DS_I[3]
  PIN IE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0024 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 157.152174 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 45.24 79.84 45.4 80 ;
    END
  END IE_I
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52976 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 140.434783 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 13.52 79.84 13.68 80 ;
    END
  END ODN_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53088 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.723602 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 11.18 79.84 11.34 80 ;
    END
  END ODP_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.78736 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.495015 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.56 79.84 14.72 80 ;
    END
  END OE_I
  PIN PD_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.996 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 156.704969 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.18 79.84 37.34 80 ;
    END
  END PD_I
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN PU_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99376 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 156.611801 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 34.32 79.84 34.48 80 ;
    END
  END PU_I
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53232 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.754658 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 22.1 79.84 22.26 80 ;
    END
  END SR_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN STE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0088 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 157.313665 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.82 79.84 40.98 80 ;
    END
  END STE_I[0]
  PIN STE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99552 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 156.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 30.68 79.84 30.84 80 ;
    END
  END STE_I[1]
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06 LAYER BA ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 0 39.576 60 40.825 ;
    END
  END VBIAS
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER YZ ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER WT ;
      RECT 0 0 60 80 ;
    LAYER BA ;
      RECT 0 0 60 80 ;
    LAYER WA ;
      RECT 0 0 60 80 ;
    LAYER BB ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_GPIO_RVT28_V

MACRO RIIO_EG1D80V_GPI_PD_RVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPI_PD_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 400.1975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 135.895 LAYER BB ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER IA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 241.9675 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 15.4548 LAYER WA ;
    ANTENNAPARTIALCUTAREA 10.4976 LAYER WT ;
    ANTENNAPARTIALCUTAREA 13.226976 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A2 ;
    ANTENNADIFFAREA 163.4 LAYER BA ;
    ANTENNADIFFAREA 163.4 LAYER C3 ;
    ANTENNADIFFAREA 163.4 LAYER BB ;
    ANTENNADIFFAREA 163.4 LAYER IA ;
    ANTENNADIFFAREA 163.4 LAYER OI ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN DI_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.02096 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.78 79.84 39.94 80 ;
    END
  END DI_O[0]
  PIN DI_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.01968 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.96 79.84 38.12 80 ;
    END
  END DI_O[1]
  PIN IE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0024 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 157.152174 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 45.24 79.84 45.4 80 ;
    END
  END IE_I
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN STE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0088 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 157.313665 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.82 79.84 40.98 80 ;
    END
  END STE_I[0]
  PIN STE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99552 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 156.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 30.68 79.84 30.84 80 ;
    END
  END STE_I[1]
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER YZ ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER WT ;
      RECT 0 0 60 80 ;
    LAYER BA ;
      RECT 0 0 60 80 ;
    LAYER WA ;
      RECT 0 0 60 80 ;
    LAYER BB ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_GPI_PD_RVT28_V

MACRO RIIO_EG1D80V_GPI_PU_RVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPI_PU_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 400.1975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 135.895 LAYER BB ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER IA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 241.9675 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 15.4548 LAYER WA ;
    ANTENNAPARTIALCUTAREA 10.4976 LAYER WT ;
    ANTENNAPARTIALCUTAREA 13.226976 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A2 ;
    ANTENNADIFFAREA 163.4 LAYER BA ;
    ANTENNADIFFAREA 163.4 LAYER C3 ;
    ANTENNADIFFAREA 163.4 LAYER BB ;
    ANTENNADIFFAREA 163.4 LAYER IA ;
    ANTENNADIFFAREA 163.4 LAYER OI ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN DI_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.02096 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.78 79.84 39.94 80 ;
    END
  END DI_O[0]
  PIN DI_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.01968 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.96 79.84 38.12 80 ;
    END
  END DI_O[1]
  PIN IE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0024 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 157.152174 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 45.24 79.84 45.4 80 ;
    END
  END IE_I
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN STE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0088 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 157.313665 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.82 79.84 40.98 80 ;
    END
  END STE_I[0]
  PIN STE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99552 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 156.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 30.68 79.84 30.84 80 ;
    END
  END STE_I[1]
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER YZ ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER WT ;
      RECT 0 0 60 80 ;
    LAYER BA ;
      RECT 0 0 60 80 ;
    LAYER WA ;
      RECT 0 0 60 80 ;
    LAYER BB ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_GPI_PU_RVT28_V

MACRO RIIO_EG1D80V_GPI_RVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPI_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 400.1975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 135.895 LAYER BB ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER IA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 241.9675 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 15.4548 LAYER WA ;
    ANTENNAPARTIALCUTAREA 10.4976 LAYER WT ;
    ANTENNAPARTIALCUTAREA 13.226976 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A2 ;
    ANTENNADIFFAREA 163.4 LAYER BA ;
    ANTENNADIFFAREA 163.4 LAYER C3 ;
    ANTENNADIFFAREA 163.4 LAYER BB ;
    ANTENNADIFFAREA 163.4 LAYER IA ;
    ANTENNADIFFAREA 163.4 LAYER OI ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN DI_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.02096 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 39.78 79.84 39.94 80 ;
    END
  END DI_O[0]
  PIN DI_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.01968 LAYER C1 ;
    ANTENNADIFFAREA 0.04048 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.96 79.84 38.12 80 ;
    END
  END DI_O[1]
  PIN IE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0024 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 157.152174 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 45.24 79.84 45.4 80 ;
    END
  END IE_I
  PIN PD_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.996 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 156.704969 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 37.18 79.84 37.34 80 ;
    END
  END PD_I
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN PU_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99376 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 156.611801 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 34.32 79.84 34.48 80 ;
    END
  END PU_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN STE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0088 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 157.313665 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 40.82 79.84 40.98 80 ;
    END
  END STE_I[0]
  PIN STE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.99552 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 156.791925 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 30.68 79.84 30.84 80 ;
    END
  END STE_I[1]
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER YZ ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER WT ;
      RECT 0 0 60 80 ;
    LAYER BA ;
      RECT 0 0 60 80 ;
    LAYER WA ;
      RECT 0 0 60 80 ;
    LAYER BB ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_GPI_RVT28_V

MACRO RIIO_EG1D80V_GPO_RVT28_V
  CLASS PAD OUTPUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPO_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52912 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.704969 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.24 79.84 19.4 80 ;
    END
  END CO_I
  PIN PAD_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 400.1975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 135.895 LAYER BB ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER IA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 241.9675 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 15.4548 LAYER WA ;
    ANTENNAPARTIALCUTAREA 10.4976 LAYER WT ;
    ANTENNAPARTIALCUTAREA 13.226976 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A2 ;
    ANTENNADIFFAREA 208.5584 LAYER BA ;
    ANTENNADIFFAREA 208.5584 LAYER C3 ;
    ANTENNADIFFAREA 208.5584 LAYER BB ;
    ANTENNADIFFAREA 208.5584 LAYER IA ;
    ANTENNADIFFAREA 208.5584 LAYER OI ;
    ANTENNADIFFAREA 208.5584 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.76592 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.287798 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 8.32 79.84 8.48 80 ;
    END
  END DO_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7984 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.962733 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 24.18 79.84 24.34 80 ;
    END
  END DS_I[0]
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.796 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.829193 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 26.78 79.84 26.94 80 ;
    END
  END DS_I[1]
  PIN DS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53232 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 140.512422 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 9.62 79.84 9.78 80 ;
    END
  END DS_I[2]
  PIN DS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52864 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.773292 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 3.9 79.84 4.06 80 ;
    END
  END DS_I[3]
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52976 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 140.434783 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 13.52 79.84 13.68 80 ;
    END
  END ODN_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53088 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.723602 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 11.18 79.84 11.34 80 ;
    END
  END ODP_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.78736 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.495015 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.56 79.84 14.72 80 ;
    END
  END OE_I
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06 LAYER BA ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 0 39.576 60 40.825 ;
    END
  END VBIAS
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53232 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.754658 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 22.1 79.84 22.26 80 ;
    END
  END SR_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER YZ ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER WT ;
      RECT 0 0 60 80 ;
    LAYER BA ;
      RECT 0 0 60 80 ;
    LAYER WA ;
      RECT 0 0 60 80 ;
    LAYER BB ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_GPO_RVT28_V

MACRO RIIO_EG1D80V_GPO_X040_RVT28_V
  CLASS PAD OUTPUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPO_X040_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52912 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.704969 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.24 79.84 19.4 80 ;
    END
  END CO_I
  PIN PAD_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 400.1975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 135.895 LAYER BB ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER IA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 241.9675 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 15.4548 LAYER WA ;
    ANTENNAPARTIALCUTAREA 10.4976 LAYER WT ;
    ANTENNAPARTIALCUTAREA 13.226976 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A2 ;
    ANTENNADIFFAREA 174.6896 LAYER BA ;
    ANTENNADIFFAREA 174.6896 LAYER C3 ;
    ANTENNADIFFAREA 174.6896 LAYER BB ;
    ANTENNADIFFAREA 174.6896 LAYER IA ;
    ANTENNADIFFAREA 174.6896 LAYER OI ;
    ANTENNADIFFAREA 174.6896 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.76592 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.287798 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 8.32 79.84 8.48 80 ;
    END
  END DO_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7984 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.959627 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 24.18 79.84 24.34 80 ;
    END
  END DS_I[0]
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.796 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.829193 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 26.78 79.84 26.94 80 ;
    END
  END DS_I[1]
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06 LAYER BA ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 0 39.576 60 40.825 ;
    END
  END VBIAS
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52976 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 140.434783 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 13.52 79.84 13.68 80 ;
    END
  END ODN_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53088 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.723602 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 11.18 79.84 11.34 80 ;
    END
  END ODP_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.78736 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.495015 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.56 79.84 14.72 80 ;
    END
  END OE_I
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53232 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.754658 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 22.1 79.84 22.26 80 ;
    END
  END SR_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER YZ ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER WT ;
      RECT 0 0 60 80 ;
    LAYER BA ;
      RECT 0 0 60 80 ;
    LAYER WA ;
      RECT 0 0 60 80 ;
    LAYER BB ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_GPO_X040_RVT28_V

MACRO RIIO_EG1D80V_GPO_X080_RVT28_V
  CLASS PAD OUTPUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPO_X080_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52912 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.704969 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.24 79.84 19.4 80 ;
    END
  END CO_I
  PIN PAD_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 400.1975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 135.895 LAYER BB ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER IA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 241.9675 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 15.4548 LAYER WA ;
    ANTENNAPARTIALCUTAREA 10.4976 LAYER WT ;
    ANTENNAPARTIALCUTAREA 13.226976 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A2 ;
    ANTENNADIFFAREA 185.9792 LAYER BA ;
    ANTENNADIFFAREA 185.9792 LAYER C3 ;
    ANTENNADIFFAREA 185.9792 LAYER BB ;
    ANTENNADIFFAREA 185.9792 LAYER IA ;
    ANTENNADIFFAREA 185.9792 LAYER OI ;
    ANTENNADIFFAREA 185.9792 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.76592 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.287798 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 8.32 79.84 8.48 80 ;
    END
  END DO_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7984 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.962733 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 24.18 79.84 24.34 80 ;
    END
  END DS_I[0]
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.796 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.829193 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 26.78 79.84 26.94 80 ;
    END
  END DS_I[1]
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06 LAYER BA ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 0 39.576 60 40.825 ;
    END
  END VBIAS
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52976 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 140.434783 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 13.52 79.84 13.68 80 ;
    END
  END ODN_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53088 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.723602 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 11.18 79.84 11.34 80 ;
    END
  END ODP_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.78736 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.495015 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.56 79.84 14.72 80 ;
    END
  END OE_I
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53232 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.754658 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 22.1 79.84 22.26 80 ;
    END
  END SR_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER YZ ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER WT ;
      RECT 0 0 60 80 ;
    LAYER BA ;
      RECT 0 0 60 80 ;
    LAYER WA ;
      RECT 0 0 60 80 ;
    LAYER BB ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_GPO_X080_RVT28_V

MACRO RIIO_EG1D80V_GPO_X120_RVT28_V
  CLASS PAD OUTPUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPO_X120_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52912 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.704969 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.24 79.84 19.4 80 ;
    END
  END CO_I
  PIN PAD_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 400.1975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 135.895 LAYER BB ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER IA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 241.9675 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 15.4548 LAYER WA ;
    ANTENNAPARTIALCUTAREA 10.4976 LAYER WT ;
    ANTENNAPARTIALCUTAREA 13.226976 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A2 ;
    ANTENNADIFFAREA 197.2688 LAYER BA ;
    ANTENNADIFFAREA 197.2688 LAYER C3 ;
    ANTENNADIFFAREA 197.2688 LAYER BB ;
    ANTENNADIFFAREA 197.2688 LAYER IA ;
    ANTENNADIFFAREA 197.2688 LAYER OI ;
    ANTENNADIFFAREA 197.2688 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.76592 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.287798 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 8.32 79.84 8.48 80 ;
    END
  END DO_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7984 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.962733 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 24.18 79.84 24.34 80 ;
    END
  END DS_I[0]
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.796 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.829193 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 26.78 79.84 26.94 80 ;
    END
  END DS_I[1]
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06 LAYER BA ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 0 39.576 60 40.825 ;
    END
  END VBIAS
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52976 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 140.434783 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 13.52 79.84 13.68 80 ;
    END
  END ODN_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53088 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.723602 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 11.18 79.84 11.34 80 ;
    END
  END ODP_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.78736 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.495015 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.56 79.84 14.72 80 ;
    END
  END OE_I
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53232 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.754658 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 22.1 79.84 22.26 80 ;
    END
  END SR_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER YZ ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER WT ;
      RECT 0 0 60 80 ;
    LAYER BA ;
      RECT 0 0 60 80 ;
    LAYER WA ;
      RECT 0 0 60 80 ;
    LAYER BB ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_GPO_X120_RVT28_V

MACRO RIIO_EG1D80V_GPO_X160_RVT28_V
  CLASS PAD OUTPUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPO_X160_RVT28_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52912 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.704969 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 19.24 79.84 19.4 80 ;
    END
  END CO_I
  PIN PAD_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 400.1975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 135.895 LAYER BB ;
    ANTENNAPARTIALMETALAREA 127.08 LAYER IA ;
    ANTENNAPARTIALMETALAREA 518.645 LAYER OI ;
    ANTENNAPARTIALMETALAREA 241.9675 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 15.4548 LAYER WA ;
    ANTENNAPARTIALCUTAREA 10.4976 LAYER WT ;
    ANTENNAPARTIALCUTAREA 13.226976 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 15.116544 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A2 ;
    ANTENNADIFFAREA 208.5584 LAYER BA ;
    ANTENNADIFFAREA 208.5584 LAYER C3 ;
    ANTENNADIFFAREA 208.5584 LAYER BB ;
    ANTENNADIFFAREA 208.5584 LAYER IA ;
    ANTENNADIFFAREA 208.5584 LAYER OI ;
    ANTENNADIFFAREA 208.5584 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER OI ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 25.35 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 25.35 ;
        RECT 30.55 0 34.15 25.35 ;
        RECT 25.85 0 29.45 25.35 ;
        RECT 21.15 0 24.75 25.35 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 25.35 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER BB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.76592 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.287798 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 8.32 79.84 8.48 80 ;
    END
  END DO_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7984 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.962733 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 24.18 79.84 24.34 80 ;
    END
  END DS_I[0]
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.796 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 187.829193 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 26.78 79.84 26.94 80 ;
    END
  END DS_I[1]
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06 LAYER BA ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 0 39.576 60 40.825 ;
    END
  END VBIAS
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.52976 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 140.434783 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 13.52 79.84 13.68 80 ;
    END
  END ODN_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53088 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.723602 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 11.18 79.84 11.34 80 ;
    END
  END ODP_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.78736 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C1 ;
      ANTENNAMAXAREACAR 18.495015 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 14.56 79.84 14.72 80 ;
    END
  END OE_I
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER OI ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER OI ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER OI ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER OI ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER OI ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER OI ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER OI ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER OI ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER OI ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER OI ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER OI ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER OI ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.53232 LAYER C1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C1 ;
      ANTENNAMAXAREACAR 138.754658 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 22.1 79.84 22.26 80 ;
    END
  END SR_I
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER YZ ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER OI ;
      RECT 0 0 60 80 ;
    LAYER JQ ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER WT ;
      RECT 0 0 60 80 ;
    LAYER BA ;
      RECT 0 0 60 80 ;
    LAYER WA ;
      RECT 0 0 60 80 ;
    LAYER BB ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_GPO_X160_RVT28_V

MACRO RIIO_EG1D80V_POR_CORE_V0D3_RVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_POR_CORE_V0D3_RVT28_V 0 0 ;
  SIZE 8 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 8 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 8 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 8 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 8 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 8 20.65 ;
    END
    PORT
      LAYER C2 ;
        RECT 0 3.325 8 5.825 ;
      LAYER IA ;
        RECT 0 3.67 8 6.55 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 0 59.35 8 62.95 ;
    END
    PORT
      LAYER C2 ;
        RECT 0 74.575 8 77.075 ;
      LAYER IA ;
        RECT 0 73.45 8 77.05 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 0 64.05 8 67.65 ;
    END
    PORT
      LAYER C2 ;
        RECT 0 70.825 8 73.325 ;
      LAYER IA ;
        RECT 0 68.75 8 72.35 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 8 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 8 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 8 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 8 15.95 ;
    END
    PORT
      LAYER C2 ;
        RECT 0 7.075 8 9.575 ;
      LAYER IA ;
        RECT 0 7.65 8 11.25 ;
    END
  END VDDIO
  PIN POR_N_CORE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8644 LAYER C1 ;
    ANTENNADIFFAREA 0.04224 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.778 79.86 5.918 80 ;
    END
  END POR_N_CORE_O
  PIN VSS_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_por VSS_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 4.998 70.825 5.138 80 ;
    END
  END VSS_POR
  PIN VDD_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd_por VDD_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 4.218 70.825 4.358 80 ;
    END
  END VDD_POR
  OBS
    LAYER CA ;
      RECT 0 0 8 80 ;
    LAYER M1 ;
      RECT 0 0 8 80 ;
    LAYER V1 ;
      RECT 0 0 8 80 ;
    LAYER M2 ;
      RECT 0 0 8 80 ;
    LAYER A1 ;
      RECT 0 0 8 80 ;
    LAYER C2 ;
      RECT 0 0 8 80 ;
    LAYER IA ;
      RECT 0 0 8 80 ;
    LAYER YZ ;
      RECT 0 0 8 80 ;
    LAYER CB ;
      RECT 0 0 8 80 ;
    LAYER OI ;
      RECT 0 0 8 80 ;
    LAYER JQ ;
      RECT 0 0 8 80 ;
    LAYER AY ;
      RECT 0 0 8 80 ;
    LAYER C1 ;
      RECT 0 0 8 80 ;
    LAYER WT ;
      RECT 0 0 8 80 ;
    LAYER BA ;
      RECT 0 0 8 80 ;
    LAYER WA ;
      RECT 0 0 8 80 ;
    LAYER BB ;
      RECT 0 0 8 80 ;
    LAYER C3 ;
      RECT 0 0 8 80 ;
    LAYER A2 ;
      RECT 0 0 8 80 ;
  END
END RIIO_EG1D80V_POR_CORE_V0D3_RVT28_V

MACRO RIIO_EG1D80V_POR_CORE_V0D5_RVT28_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_POR_CORE_V0D5_RVT28_V 0 0 ;
  SIZE 8 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 0 54.65 8 58.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 45.25 8 48.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 40.55 8 44.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 26.45 8 30.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 17.05 8 20.65 ;
    END
    PORT
      LAYER C2 ;
        RECT 0 3.325 8 5.825 ;
      LAYER IA ;
        RECT 0 3.67 8 6.55 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 0 59.35 8 62.95 ;
    END
    PORT
      LAYER C2 ;
        RECT 0 74.575 8 77.075 ;
      LAYER IA ;
        RECT 0 73.45 8 77.05 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 0 64.05 8 67.65 ;
    END
    PORT
      LAYER C2 ;
        RECT 0 70.825 8 73.325 ;
      LAYER IA ;
        RECT 0 68.75 8 72.35 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 0 49.95 8 53.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.85 8 39.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 31.15 8 34.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 12.35 8 15.95 ;
    END
    PORT
      LAYER C2 ;
        RECT 0 7.075 8 9.575 ;
      LAYER IA ;
        RECT 0 7.65 8 11.25 ;
    END
  END VDDIO
  PIN POR_N_CORE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9344 LAYER C1 ;
    ANTENNADIFFAREA 0.04224 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 5.778 79.86 5.918 80 ;
    END
  END POR_N_CORE_O
  PIN VSS_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_por VSS_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 4.998 70.825 5.138 80 ;
    END
  END VSS_POR
  PIN VDD_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd_por VDD_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 4.218 70.825 4.358 80 ;
    END
  END VDD_POR
  OBS
    LAYER CA ;
      RECT 0 0 8 80 ;
    LAYER M1 ;
      RECT 0 0 8 80 ;
    LAYER V1 ;
      RECT 0 0 8 80 ;
    LAYER M2 ;
      RECT 0 0 8 80 ;
    LAYER A1 ;
      RECT 0 0 8 80 ;
    LAYER C2 ;
      RECT 0 0 8 80 ;
    LAYER IA ;
      RECT 0 0 8 80 ;
    LAYER YZ ;
      RECT 0 0 8 80 ;
    LAYER CB ;
      RECT 0 0 8 80 ;
    LAYER OI ;
      RECT 0 0 8 80 ;
    LAYER JQ ;
      RECT 0 0 8 80 ;
    LAYER AY ;
      RECT 0 0 8 80 ;
    LAYER C1 ;
      RECT 0 0 8 80 ;
    LAYER WT ;
      RECT 0 0 8 80 ;
    LAYER BA ;
      RECT 0 0 8 80 ;
    LAYER WA ;
      RECT 0 0 8 80 ;
    LAYER BB ;
      RECT 0 0 8 80 ;
    LAYER C3 ;
      RECT 0 0 8 80 ;
    LAYER A2 ;
      RECT 0 0 8 80 ;
  END
END RIIO_EG1D80V_POR_CORE_V0D5_RVT28_V

MACRO RIIO_EG1D80V_BIAS_RVT28_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_BIAS_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER OI ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER OI ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER OI ;
        RECT 0 2.35 58.25 5.95 ;
        RECT 0 11.75 58.25 15.35 ;
        RECT 0 44.65 58.25 48.25 ;
        RECT 0 54.05 58.25 57.65 ;
        RECT 0 21.15 58.249 24.75 ;
        RECT 0 35.25 58.249 38.85 ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 49.35 25.35 52.95 ;
      LAYER IA ;
        RECT 54.65 0 58.25 60 ;
        RECT 45.25 0 48.85 60 ;
        RECT 40.55 0 44.15 60 ;
        RECT 26.45 0 30.05 60 ;
        RECT 17.05 0 20.65 60 ;
        RECT 3.67 0 6.55 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.352 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 39.575 0 40.825 60 ;
    END
  END VBIAS
  PIN VTMP_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9 LAYER C2 ;
    ANTENNADIFFAREA 0.32 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.4 LAYER C2 ;
      ANTENNAMAXAREACAR 1.783129 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.935 80 28.095 ;
    END
  END VTMP_O
  PIN VBG_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9 LAYER C2 ;
    ANTENNADIFFAREA 0.32 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.4 LAYER C2 ;
      ANTENNAMAXAREACAR 2.083058 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.115 80 26.275 ;
    END
  END VBG_O
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN TRIM_VBG_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7496 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03808 LAYER C2 ;
      ANTENNAMAXAREACAR 301.585003 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 40.26 80 40.42 ;
    END
  END TRIM_VBG_I[4]
  PIN TRIM_VBG_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7496 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03808 LAYER C2 ;
      ANTENNAMAXAREACAR 301.070297 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 40 80 40.16 ;
    END
  END TRIM_VBG_I[3]
  PIN TRIM_VBG_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7496 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04704 LAYER C2 ;
      ANTENNAMAXAREACAR 251.095557 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 39.74 80 39.9 ;
    END
  END TRIM_VBG_I[2]
  PIN TRIM_VBG_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7496 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.07392 LAYER C2 ;
      ANTENNAMAXAREACAR 165.619755 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 39.48 80 39.64 ;
    END
  END TRIM_VBG_I[1]
  PIN TRIM_VBG_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7496 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1456 LAYER C2 ;
      ANTENNAMAXAREACAR 85.576374 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 39.22 80 39.38 ;
    END
  END TRIM_VBG_I[0]
  PIN TRIM_CURV_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7496 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03808 LAYER C2 ;
      ANTENNAMAXAREACAR 299.192469 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 42.34 80 42.5 ;
    END
  END TRIM_CURV_I[4]
  PIN TRIM_CURV_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7496 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03808 LAYER C2 ;
      ANTENNAMAXAREACAR 298.129121 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 42.08 80 42.24 ;
    END
  END TRIM_CURV_I[3]
  PIN TRIM_CURV_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7496 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04704 LAYER C2 ;
      ANTENNAMAXAREACAR 246.496599 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 41.82 80 41.98 ;
    END
  END TRIM_CURV_I[2]
  PIN TRIM_CURV_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7496 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.07392 LAYER C2 ;
      ANTENNAMAXAREACAR 162.755073 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 41.56 80 41.72 ;
    END
  END TRIM_CURV_I[1]
  PIN TRIM_CURV_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7496 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1456 LAYER C2 ;
      ANTENNAMAXAREACAR 84.333516 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 41.3 80 41.46 ;
    END
  END TRIM_CURV_I[0]
  PIN TRIM_BIAS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 214.284161 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 48.28 80 48.44 ;
    END
  END TRIM_BIAS_I[3]
  PIN TRIM_BIAS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8984 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 191.787267 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 47.76 80 47.92 ;
    END
  END TRIM_BIAS_I[2]
  PIN TRIM_BIAS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7336 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 146.43323 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 47.24 80 47.4 ;
    END
  END TRIM_BIAS_I[1]
  PIN TRIM_BIAS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.316 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 169.290373 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 46.72 80 46.88 ;
    END
  END TRIM_BIAS_I[0]
  PIN IBIAS_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 24.815 80 24.975 ;
    END
  END IBIAS_O[9]
  PIN IBIAS_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 24.555 80 24.715 ;
    END
  END IBIAS_O[8]
  PIN IBIAS_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 23.255 80 23.415 ;
    END
  END IBIAS_O[7]
  PIN IBIAS_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 22.995 80 23.155 ;
    END
  END IBIAS_O[6]
  PIN IBIAS_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 22.735 80 22.895 ;
    END
  END IBIAS_O[5]
  PIN IBIAS_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 22.475 80 22.635 ;
    END
  END IBIAS_O[4]
  PIN IBIAS_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 21.695 80 21.855 ;
    END
  END IBIAS_O[3]
  PIN IBIAS_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 21.435 80 21.595 ;
    END
  END IBIAS_O[2]
  PIN IBIAS_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 21.175 80 21.335 ;
    END
  END IBIAS_O[1]
  PIN IBIAS_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.415 80 27.575 ;
    END
  END IBIAS_O[15]
  PIN IBIAS_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.155 80 27.315 ;
    END
  END IBIAS_O[14]
  PIN IBIAS_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.895 80 27.055 ;
    END
  END IBIAS_O[13]
  PIN IBIAS_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.635 80 26.795 ;
    END
  END IBIAS_O[12]
  PIN EN_VBIAS_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5688 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 101.439441 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 50.62 80 50.78 ;
    END
  END EN_VBIAS_I
  PIN IBIAS_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 20.915 80 21.075 ;
    END
  END IBIAS_O[0]
  PIN IBIAS_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 25.075 80 25.235 ;
    END
  END IBIAS_O[10]
  PIN IBIAS_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6936 LAYER C2 ;
    ANTENNADIFFAREA 0.088 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 25.335 80 25.495 ;
    END
  END IBIAS_O[11]
  PIN EN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1512 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 123.936335 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 50.1 80 50.26 ;
    END
  END EN_I
  PIN BG_STARTUP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6488 LAYER C2 ;
    ANTENNADIFFAREA 0.2528 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.474 LAYER C2 ;
      ANTENNAMAXAREACAR 9.520777 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 49.58 80 49.74 ;
    END
  END BG_STARTUP_I
  PIN BG_VALID_N_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9816 LAYER C2 ;
    ANTENNADIFFAREA 0.1045 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.099 LAYER C2 ;
      ANTENNAMAXAREACAR 21.908232 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 49.06 80 49.22 ;
    END
  END BG_VALID_N_O
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER YZ ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER WT ;
      RECT 0 0 80 60 ;
    LAYER BA ;
      RECT 0 0 80 60 ;
    LAYER WA ;
      RECT 0 0 80 60 ;
    LAYER BB ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_BIAS_RVT28_H

MACRO RIIO_EG1D80V_GPIO_RVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPIO_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.555 LAYER BB ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER IA ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER OI ;
    ANTENNAPARTIALMETALAREA 33.7006 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 16.2324 LAYER WA ;
    ANTENNAPARTIALCUTAREA 19.8288 LAYER WT ;
    ANTENNAPARTIALCUTAREA 12.387168 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.4472 LAYER A2 ;
    ANTENNADIFFAREA 193.746 LAYER BA ;
    ANTENNADIFFAREA 193.746 LAYER C3 ;
    ANTENNADIFFAREA 193.746 LAYER BB ;
    ANTENNADIFFAREA 193.746 LAYER IA ;
    ANTENNADIFFAREA 193.746 LAYER OI ;
    ANTENNADIFFAREA 193.746 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BB ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.26208 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 132.226708 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.06 80 27.22 ;
    END
  END CO_I
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.67808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 146.583851 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.58 80 27.74 ;
    END
  END SR_I
  PIN DI_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.55648 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 29.66 80 29.82 ;
    END
  END DI_O[0]
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.59808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 8.623363 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.4 80 3.56 ;
    END
  END OE_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.82368 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 44.208075 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.02 80 26.18 ;
    END
  END ODP_I
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51504 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 67.431677 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.54 80 26.7 ;
    END
  END ODN_I
  PIN IE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.80768 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 46.139752 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 29.14 80 29.3 ;
    END
  END IE_I
  PIN STE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.09568 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 124.018634 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 31.22 80 31.38 ;
    END
  END STE_I[1]
  PIN PD_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.09728 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 99.630435 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 28.62 80 28.78 ;
    END
  END PD_I
  PIN PU_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.55488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 120.456522 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 28.1 80 28.26 ;
    END
  END PU_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.88608 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 213.965839 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 23.94 80 24.1 ;
    END
  END DS_I[0]
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.55488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 13.466369 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.92 80 4.08 ;
    END
  END DO_I
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 39.575 0 40.825 60 ;
    END
  END VBIAS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.42688 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 192.76087 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 24.46 80 24.62 ;
    END
  END DS_I[1]
  PIN DS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.55488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 116.860248 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 24.98 80 25.14 ;
    END
  END DS_I[2]
  PIN DS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.09728 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 95.86646 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 25.5 80 25.66 ;
    END
  END DS_I[3]
  PIN STE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 65.021739 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 30.7 80 30.86 ;
    END
  END STE_I[0]
  PIN DI_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.85008 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 30.18 80 30.34 ;
    END
  END DI_O[1]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER YZ ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER WT ;
      RECT 0 0 80 60 ;
    LAYER BA ;
      RECT 0 0 80 60 ;
    LAYER WA ;
      RECT 0 0 80 60 ;
    LAYER BB ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_GPIO_RVT28_H

MACRO RIIO_EG1D80V_GPI_PD_RVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPI_PD_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.555 LAYER BB ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER IA ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER OI ;
    ANTENNAPARTIALMETALAREA 33.7006 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 16.2324 LAYER WA ;
    ANTENNAPARTIALCUTAREA 19.8288 LAYER WT ;
    ANTENNAPARTIALCUTAREA 12.387168 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.4472 LAYER A2 ;
    ANTENNADIFFAREA 148.5876 LAYER BA ;
    ANTENNADIFFAREA 148.5876 LAYER C3 ;
    ANTENNADIFFAREA 148.5876 LAYER BB ;
    ANTENNADIFFAREA 148.5876 LAYER IA ;
    ANTENNADIFFAREA 148.5876 LAYER OI ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BB ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN DI_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.55648 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 29.66 80 29.82 ;
    END
  END DI_O[0]
  PIN IE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.80768 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 46.139752 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 29.14 80 29.3 ;
    END
  END IE_I
  PIN STE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.09568 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 124.018634 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 31.22 80 31.38 ;
    END
  END STE_I[1]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN STE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 65.021739 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 30.7 80 30.86 ;
    END
  END STE_I[0]
  PIN DI_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.85008 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 30.18 80 30.34 ;
    END
  END DI_O[1]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER YZ ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER WT ;
      RECT 0 0 80 60 ;
    LAYER BA ;
      RECT 0 0 80 60 ;
    LAYER WA ;
      RECT 0 0 80 60 ;
    LAYER BB ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_GPI_PD_RVT28_H

MACRO RIIO_EG1D80V_GPI_PU_RVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPI_PU_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.555 LAYER BB ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER IA ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER OI ;
    ANTENNAPARTIALMETALAREA 33.7006 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 16.2324 LAYER WA ;
    ANTENNAPARTIALCUTAREA 19.8288 LAYER WT ;
    ANTENNAPARTIALCUTAREA 12.387168 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.4472 LAYER A2 ;
    ANTENNADIFFAREA 148.5876 LAYER BA ;
    ANTENNADIFFAREA 148.5876 LAYER C3 ;
    ANTENNADIFFAREA 148.5876 LAYER BB ;
    ANTENNADIFFAREA 148.5876 LAYER IA ;
    ANTENNADIFFAREA 148.5876 LAYER OI ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BB ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN DI_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.55648 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 29.66 80 29.82 ;
    END
  END DI_O[0]
  PIN IE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.80768 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 46.139752 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 29.14 80 29.3 ;
    END
  END IE_I
  PIN STE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.09568 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 124.018634 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 31.22 80 31.38 ;
    END
  END STE_I[1]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN STE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 65.021739 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 30.7 80 30.86 ;
    END
  END STE_I[0]
  PIN DI_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.85008 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 30.18 80 30.34 ;
    END
  END DI_O[1]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER YZ ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER WT ;
      RECT 0 0 80 60 ;
    LAYER BA ;
      RECT 0 0 80 60 ;
    LAYER WA ;
      RECT 0 0 80 60 ;
    LAYER BB ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_GPI_PU_RVT28_H

MACRO RIIO_EG1D80V_GPI_RVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPI_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.555 LAYER BB ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER IA ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER OI ;
    ANTENNAPARTIALMETALAREA 33.7006 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 16.2324 LAYER WA ;
    ANTENNAPARTIALCUTAREA 19.8288 LAYER WT ;
    ANTENNAPARTIALCUTAREA 12.387168 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.4472 LAYER A2 ;
    ANTENNADIFFAREA 148.5876 LAYER BA ;
    ANTENNADIFFAREA 148.5876 LAYER C3 ;
    ANTENNADIFFAREA 148.5876 LAYER BB ;
    ANTENNADIFFAREA 148.5876 LAYER IA ;
    ANTENNADIFFAREA 148.5876 LAYER OI ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BB ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN DI_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.55648 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 29.66 80 29.82 ;
    END
  END DI_O[0]
  PIN IE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.80768 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 46.139752 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 29.14 80 29.3 ;
    END
  END IE_I
  PIN STE_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.09568 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 124.018634 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 31.22 80 31.38 ;
    END
  END STE_I[1]
  PIN PD_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.09728 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 99.630435 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 28.62 80 28.78 ;
    END
  END PD_I
  PIN PU_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.55488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 120.456522 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 28.1 80 28.26 ;
    END
  END PU_I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN STE_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 65.021739 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 30.7 80 30.86 ;
    END
  END STE_I[0]
  PIN DI_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.85008 LAYER C2 ;
    ANTENNADIFFAREA 0.04048 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 30.18 80 30.34 ;
    END
  END DI_O[1]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER YZ ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER WT ;
      RECT 0 0 80 60 ;
    LAYER BA ;
      RECT 0 0 80 60 ;
    LAYER WA ;
      RECT 0 0 80 60 ;
    LAYER BB ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_GPI_RVT28_H

MACRO RIIO_EG1D80V_GPO_RVT28_H
  CLASS PAD OUTPUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPO_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN PAD_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.555 LAYER BB ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER IA ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER OI ;
    ANTENNAPARTIALMETALAREA 33.7006 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 16.2324 LAYER WA ;
    ANTENNAPARTIALCUTAREA 19.8288 LAYER WT ;
    ANTENNAPARTIALCUTAREA 12.387168 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.4472 LAYER A2 ;
    ANTENNADIFFAREA 193.746 LAYER BA ;
    ANTENNADIFFAREA 193.746 LAYER C3 ;
    ANTENNADIFFAREA 193.746 LAYER BB ;
    ANTENNADIFFAREA 193.746 LAYER IA ;
    ANTENNADIFFAREA 193.746 LAYER OI ;
    ANTENNADIFFAREA 193.746 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BB ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.26208 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 132.226708 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.06 80 27.22 ;
    END
  END CO_I
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.67808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 146.583851 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.58 80 27.74 ;
    END
  END SR_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.59808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 8.623363 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.4 80 3.56 ;
    END
  END OE_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.82368 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 44.208075 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.02 80 26.18 ;
    END
  END ODP_I
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51504 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 67.431677 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.54 80 26.7 ;
    END
  END ODN_I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.88608 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 213.965839 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 23.94 80 24.1 ;
    END
  END DS_I[0]
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.55488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 13.466369 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.92 80 4.08 ;
    END
  END DO_I
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 39.575 0 40.825 60 ;
    END
  END VBIAS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.42688 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 192.76087 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 24.46 80 24.62 ;
    END
  END DS_I[1]
  PIN DS_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.55488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 116.860248 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 24.98 80 25.14 ;
    END
  END DS_I[2]
  PIN DS_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.09728 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 95.86646 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 25.5 80 25.66 ;
    END
  END DS_I[3]
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER YZ ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER WT ;
      RECT 0 0 80 60 ;
    LAYER BA ;
      RECT 0 0 80 60 ;
    LAYER WA ;
      RECT 0 0 80 60 ;
    LAYER BB ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_GPO_RVT28_H

MACRO RIIO_EG1D80V_GPO_X040_RVT28_H
  CLASS PAD OUTPUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPO_X040_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN PAD_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.555 LAYER BB ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER IA ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER OI ;
    ANTENNAPARTIALMETALAREA 33.7006 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 16.2324 LAYER WA ;
    ANTENNAPARTIALCUTAREA 19.8288 LAYER WT ;
    ANTENNAPARTIALCUTAREA 12.387168 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.4472 LAYER A2 ;
    ANTENNADIFFAREA 159.8772 LAYER BA ;
    ANTENNADIFFAREA 159.8772 LAYER C3 ;
    ANTENNADIFFAREA 159.8772 LAYER BB ;
    ANTENNADIFFAREA 159.8772 LAYER IA ;
    ANTENNADIFFAREA 159.8772 LAYER OI ;
    ANTENNADIFFAREA 159.8772 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BB ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.26208 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 132.226708 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.06 80 27.22 ;
    END
  END CO_I
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.67808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 146.583851 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.58 80 27.74 ;
    END
  END SR_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.59808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 8.623363 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.4 80 3.56 ;
    END
  END OE_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.82368 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 44.208075 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.02 80 26.18 ;
    END
  END ODP_I
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51504 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 67.431677 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.54 80 26.7 ;
    END
  END ODN_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.88608 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 213.965839 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 23.94 80 24.1 ;
    END
  END DS_I[0]
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.55488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 13.466369 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.92 80 4.08 ;
    END
  END DO_I
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 39.575 0 40.825 60 ;
    END
  END VBIAS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.42688 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 192.76087 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 24.46 80 24.62 ;
    END
  END DS_I[1]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER YZ ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER WT ;
      RECT 0 0 80 60 ;
    LAYER BA ;
      RECT 0 0 80 60 ;
    LAYER WA ;
      RECT 0 0 80 60 ;
    LAYER BB ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_GPO_X040_RVT28_H

MACRO RIIO_EG1D80V_GPO_X080_RVT28_H
  CLASS PAD OUTPUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPO_X080_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN PAD_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.555 LAYER BB ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER IA ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER OI ;
    ANTENNAPARTIALMETALAREA 33.7006 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 16.2324 LAYER WA ;
    ANTENNAPARTIALCUTAREA 19.8288 LAYER WT ;
    ANTENNAPARTIALCUTAREA 12.387168 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.4472 LAYER A2 ;
    ANTENNADIFFAREA 171.1668 LAYER BA ;
    ANTENNADIFFAREA 171.1668 LAYER C3 ;
    ANTENNADIFFAREA 171.1668 LAYER BB ;
    ANTENNADIFFAREA 171.1668 LAYER IA ;
    ANTENNADIFFAREA 171.1668 LAYER OI ;
    ANTENNADIFFAREA 171.1668 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BB ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.26208 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 132.226708 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.06 80 27.22 ;
    END
  END CO_I
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.67808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 146.583851 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.58 80 27.74 ;
    END
  END SR_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.59808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 8.623363 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.4 80 3.56 ;
    END
  END OE_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.82368 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 44.208075 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.02 80 26.18 ;
    END
  END ODP_I
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51504 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 67.431677 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.54 80 26.7 ;
    END
  END ODN_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.88608 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 213.965839 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 23.94 80 24.1 ;
    END
  END DS_I[0]
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.55488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 13.466369 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.92 80 4.08 ;
    END
  END DO_I
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 39.575 0 40.825 60 ;
    END
  END VBIAS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.42688 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 192.76087 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 24.46 80 24.62 ;
    END
  END DS_I[1]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER YZ ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER WT ;
      RECT 0 0 80 60 ;
    LAYER BA ;
      RECT 0 0 80 60 ;
    LAYER WA ;
      RECT 0 0 80 60 ;
    LAYER BB ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_GPO_X080_RVT28_H

MACRO RIIO_EG1D80V_GPO_X120_RVT28_H
  CLASS PAD OUTPUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPO_X120_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN PAD_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.555 LAYER BB ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER IA ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER OI ;
    ANTENNAPARTIALMETALAREA 33.7006 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 16.2324 LAYER WA ;
    ANTENNAPARTIALCUTAREA 19.8288 LAYER WT ;
    ANTENNAPARTIALCUTAREA 12.387168 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.4472 LAYER A2 ;
    ANTENNADIFFAREA 182.4564 LAYER BA ;
    ANTENNADIFFAREA 182.4564 LAYER C3 ;
    ANTENNADIFFAREA 182.4564 LAYER BB ;
    ANTENNADIFFAREA 182.4564 LAYER IA ;
    ANTENNADIFFAREA 182.4564 LAYER OI ;
    ANTENNADIFFAREA 182.4564 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BB ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.26208 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 132.226708 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.06 80 27.22 ;
    END
  END CO_I
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.67808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 146.583851 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.58 80 27.74 ;
    END
  END SR_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.59808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 8.623363 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.4 80 3.56 ;
    END
  END OE_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.82368 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 44.208075 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.02 80 26.18 ;
    END
  END ODP_I
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51504 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 67.431677 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.54 80 26.7 ;
    END
  END ODN_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.88608 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 213.965839 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 23.94 80 24.1 ;
    END
  END DS_I[0]
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.55488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 13.466369 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.92 80 4.08 ;
    END
  END DO_I
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 39.575 0 40.825 60 ;
    END
  END VBIAS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.42688 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 192.76087 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 24.46 80 24.62 ;
    END
  END DS_I[1]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER YZ ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER WT ;
      RECT 0 0 80 60 ;
    LAYER BA ;
      RECT 0 0 80 60 ;
    LAYER WA ;
      RECT 0 0 80 60 ;
    LAYER BB ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_GPO_X120_RVT28_H

MACRO RIIO_EG1D80V_GPO_X160_RVT28_H
  CLASS PAD OUTPUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_GPO_X160_RVT28_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN PAD_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER BA ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 105.555 LAYER BB ;
    ANTENNAPARTIALMETALAREA 302.645 LAYER IA ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER OI ;
    ANTENNAPARTIALMETALAREA 33.7006 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 16.2324 LAYER WA ;
    ANTENNAPARTIALCUTAREA 19.8288 LAYER WT ;
    ANTENNAPARTIALCUTAREA 12.387168 LAYER YZ ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER JQ ;
    ANTENNAPARTIALCUTAREA 5.4472 LAYER A2 ;
    ANTENNADIFFAREA 193.746 LAYER BA ;
    ANTENNADIFFAREA 193.746 LAYER C3 ;
    ANTENNADIFFAREA 193.746 LAYER BB ;
    ANTENNADIFFAREA 193.746 LAYER IA ;
    ANTENNADIFFAREA 193.746 LAYER OI ;
    ANTENNADIFFAREA 193.746 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER BB ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER OI ;
        RECT 0 7.05 25.35 10.65 ;
        RECT 0 21.15 25.35 24.75 ;
        RECT 0 25.85 25.35 29.45 ;
        RECT 0 30.55 25.35 34.15 ;
        RECT 0 35.25 25.35 38.85 ;
        RECT 0 49.35 25.35 52.95 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN CO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.26208 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 132.226708 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.06 80 27.22 ;
    END
  END CO_I
  PIN SR_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.67808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 146.583851 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 27.58 80 27.74 ;
    END
  END SR_I
  PIN OE_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.59808 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 8.623363 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.4 80 3.56 ;
    END
  END OE_I
  PIN ODP_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.82368 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 44.208075 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.02 80 26.18 ;
    END
  END ODP_I
  PIN ODN_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51504 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 67.431677 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 26.54 80 26.7 ;
    END
  END ODN_I
  PIN DS_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.88608 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 213.965839 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 23.94 80 24.1 ;
    END
  END DS_I[0]
  PIN DO_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.55488 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21504 LAYER C2 ;
      ANTENNAMAXAREACAR 13.466369 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 3.92 80 4.08 ;
    END
  END DO_I
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER OI ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER OI ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER OI ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER OI ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER OI ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER OI ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3465 LAYER BA ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER BA ;
        RECT 39.575 0 40.825 60 ;
    END
  END VBIAS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN DS_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.42688 LAYER C2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02576 LAYER C2 ;
      ANTENNAMAXAREACAR 192.76087 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.84 24.46 80 24.62 ;
    END
  END DS_I[1]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER OI ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER OI ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER OI ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER OI ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER OI ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER OI ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER YZ ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER OI ;
      RECT 0 0 80 60 ;
    LAYER JQ ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER WT ;
      RECT 0 0 80 60 ;
    LAYER BA ;
      RECT 0 0 80 60 ;
    LAYER WA ;
      RECT 0 0 80 60 ;
    LAYER BB ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_GPO_X160_RVT28_H

MACRO RIIO_EG1D80V_POR_CORE_V0D3_RVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_POR_CORE_V0D3_RVT28_H 0 0 ;
  SIZE 80 BY 8 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 8 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 8 ;
      LAYER C3 ;
        RECT 14.573 0 17.073 8 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 8 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 8 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 8 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 8 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 8 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 8 ;
      LAYER C3 ;
        RECT 70.825 0 73.325 8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 8 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 8 ;
      LAYER C3 ;
        RECT 74.575 0 77.075 8 ;
    END
  END VSS
  PIN VSS_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_por VSS_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 70.825 2.625 80 3.125 ;
    END
  END VSS_POR
  PIN VDD_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd_por VDD_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 70.825 1.875 80 2.375 ;
    END
  END VDD_POR
  PIN POR_N_CORE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.324 LAYER C2 ;
    ANTENNADIFFAREA 0.04224 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.5 3.375 80 3.875 ;
    END
  END POR_N_CORE_O
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 8 ;
        RECT 7.65 0 11.25 8 ;
      LAYER C3 ;
        RECT 10.825 0 13.325 8 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 8 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 8 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 8 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 8 ;
    LAYER M1 ;
      RECT 0 0 80 8 ;
    LAYER V1 ;
      RECT 0 0 80 8 ;
    LAYER M2 ;
      RECT 0 0 80 8 ;
    LAYER A1 ;
      RECT 0 0 80 8 ;
    LAYER C2 ;
      RECT 0 0 80 8 ;
    LAYER IA ;
      RECT 0 0 80 8 ;
    LAYER YZ ;
      RECT 0 0 80 8 ;
    LAYER CB ;
      RECT 0 0 80 8 ;
    LAYER OI ;
      RECT 0 0 80 8 ;
    LAYER JQ ;
      RECT 0 0 80 8 ;
    LAYER AY ;
      RECT 0 0 80 8 ;
    LAYER C1 ;
      RECT 0 0 80 8 ;
    LAYER WT ;
      RECT 0 0 80 8 ;
    LAYER BA ;
      RECT 0 0 80 8 ;
    LAYER WA ;
      RECT 0 0 80 8 ;
    LAYER BB ;
      RECT 0 0 80 8 ;
    LAYER C3 ;
      RECT 0 0 80 8 ;
    LAYER A2 ;
      RECT 0 0 80 8 ;
  END
END RIIO_EG1D80V_POR_CORE_V0D3_RVT28_H

MACRO RIIO_EG1D80V_POR_CORE_V0D5_RVT28_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_POR_CORE_V0D5_RVT28_H 0 0 ;
  SIZE 80 BY 8 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IA ;
        RECT 3.67 0 6.55 8 ;
    END
    PORT
      LAYER IA ;
        RECT 17.05 0 20.65 8 ;
      LAYER C3 ;
        RECT 14.573 0 17.073 8 ;
    END
    PORT
      LAYER IA ;
        RECT 26.45 0 30.05 8 ;
    END
    PORT
      LAYER IA ;
        RECT 40.55 0 44.15 8 ;
    END
    PORT
      LAYER IA ;
        RECT 45.25 0 48.85 8 ;
    END
    PORT
      LAYER IA ;
        RECT 54.65 0 58.25 8 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IA ;
        RECT 64.05 0 67.65 8 ;
    END
    PORT
      LAYER IA ;
        RECT 68.75 0 72.35 8 ;
      LAYER C3 ;
        RECT 70.825 0 73.325 8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IA ;
        RECT 59.35 0 62.95 8 ;
    END
    PORT
      LAYER IA ;
        RECT 73.45 0 77.05 8 ;
      LAYER C3 ;
        RECT 74.575 0 77.075 8 ;
    END
  END VSS
  PIN VSS_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_por VSS_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 70.825 2.625 80 3.125 ;
    END
  END VSS_POR
  PIN VDD_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd_por VDD_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 70.825 1.875 80 2.375 ;
    END
  END VDD_POR
  PIN POR_N_CORE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.324 LAYER C2 ;
    ANTENNADIFFAREA 0.04224 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.5 3.375 80 3.875 ;
    END
  END POR_N_CORE_O
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IA ;
        RECT 12.35 0 15.95 8 ;
        RECT 7.65 0 11.25 8 ;
      LAYER C3 ;
        RECT 10.825 0 13.325 8 ;
    END
    PORT
      LAYER IA ;
        RECT 31.15 0 34.75 8 ;
    END
    PORT
      LAYER IA ;
        RECT 35.85 0 39.45 8 ;
    END
    PORT
      LAYER IA ;
        RECT 49.95 0 53.55 8 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 8 ;
    LAYER M1 ;
      RECT 0 0 80 8 ;
    LAYER V1 ;
      RECT 0 0 80 8 ;
    LAYER M2 ;
      RECT 0 0 80 8 ;
    LAYER A1 ;
      RECT 0 0 80 8 ;
    LAYER C2 ;
      RECT 0 0 80 8 ;
    LAYER IA ;
      RECT 0 0 80 8 ;
    LAYER YZ ;
      RECT 0 0 80 8 ;
    LAYER CB ;
      RECT 0 0 80 8 ;
    LAYER OI ;
      RECT 0 0 80 8 ;
    LAYER JQ ;
      RECT 0 0 80 8 ;
    LAYER AY ;
      RECT 0 0 80 8 ;
    LAYER C1 ;
      RECT 0 0 80 8 ;
    LAYER WT ;
      RECT 0 0 80 8 ;
    LAYER BA ;
      RECT 0 0 80 8 ;
    LAYER WA ;
      RECT 0 0 80 8 ;
    LAYER BB ;
      RECT 0 0 80 8 ;
    LAYER C3 ;
      RECT 0 0 80 8 ;
    LAYER A2 ;
      RECT 0 0 80 8 ;
  END
END RIIO_EG1D80V_POR_CORE_V0D5_RVT28_H

END LIBRARY
