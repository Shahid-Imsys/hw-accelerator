library ieee;
use ieee.std_logic_1164.all;
use work.all;
use work.pe1_gp_pkg.all;

entity PE_pair_top is
  generic ( USE_ASIC_MEMORIES : boolean := false );
  port (
    --Data interface --Added by CJ
    C1_REQ    : out std_logic;
    C1_REQ_RD : out std_logic;
    C2_REQ    : out std_logic;
    C2_REQ_RD : out std_logic;
    C1_ACK    : in std_logic;
    C2_ACK    : in std_logic;
    C1_REQ_D  : out std_logic_vector(159 downto 0);
    C2_REQ_D  : out std_logic_vector(159 downto 0);
    C1_IN_D   : in std_logic_vector(127 downto 0);
    C2_IN_D   : in std_logic_vector(127 downto 0);
    C1_DDI_VLD : in std_logic;
    C2_DDI_VLD : in std_logic;
    C1_RDY     : out std_logic;
    C2_RDY     : out std_logic;
    EXE        : in std_logic;
    RESUME     : in std_logic;
    C1_ID      : in std_logic_vector(5 downto 0);
    C2_ID      : in std_logic_vector(5 downto 0);


    -- clocks and control signals
    HCLK       : in    std_logic;                  -- clk input, use this or an internally generated clock for CPU core
    EVEN_C     : in    std_logic;                  -- even pulses of HCLK. Used to generate clk_e_pos and clk_e_neg.
    MRESET     : in    std_logic;                  -- system reset               low active --generated by cc
    MIRQOUT    : out   std_logic;                  -- interrupt request output
    MCKOUT1    : out   std_logic;                  -- programable clock out
    MBYPASS    : in    std_logic;
    -- SW debug
    MSDIN      : in    std_logic;                  -- serial data in (debug)
    MSDOUT     : out   std_logic;                  -- serial data out

    MLP_PWR_OK : in    std_logic;                  -- Power on indecator --From Host directly
    MWAKEUP_LP  : in    std_logic

  );
end PE_pair_top;

architecture struct of PE_pair_top is

  component SNPS_RF_SP_UHS_256x64 is
    port (
      Q        : out std_logic_vector(63 downto 0);
      ADR      : in  std_logic_vector(7 downto 0);
      D        : in  std_logic_vector(63 downto 0);
      WE       : in  std_logic;
      ME       : in  std_logic;
      CLK      : in  std_logic;
      TEST1    : in  std_logic;
      TEST_RNM : in  std_logic;
      RME      : in  std_logic;
      RM       : in  std_logic_vector(3 downto 0);
      WA       : in  std_logic_vector(1 downto 0);
      WPULSE   : in  std_logic_vector(2 downto 0);
      LS       : in  std_logic;
      BC0      : in  std_logic;
      BC1      : in  std_logic;
      BC2      : in  std_logic);
  end component;

  --RAM 0
  component FPGA_SU180_256X128X1BM1A
  port(
      A0                          :   IN   std_logic;
      A1                          :   IN   std_logic;
      A2                          :   IN   std_logic;
      A3                          :   IN   std_logic;
      A4                          :   IN   std_logic;
      A5                          :   IN   std_logic;
      A6                          :   IN   std_logic;
      A7                          :   IN   std_logic;
      DO0                         :   OUT   std_logic;
      DO1                         :   OUT   std_logic;
      DO2                         :   OUT   std_logic;
      DO3                         :   OUT   std_logic;
      DO4                         :   OUT   std_logic;
      DO5                         :   OUT   std_logic;
      DO6                         :   OUT   std_logic;
      DO7                         :   OUT   std_logic;
      DO8                         :   OUT   std_logic;
      DO9                         :   OUT   std_logic;
      DO10                        :   OUT   std_logic;
      DO11                        :   OUT   std_logic;
      DO12                        :   OUT   std_logic;
      DO13                        :   OUT   std_logic;
      DO14                        :   OUT   std_logic;
      DO15                        :   OUT   std_logic;
      DO16                        :   OUT   std_logic;
      DO17                        :   OUT   std_logic;
      DO18                        :   OUT   std_logic;
      DO19                        :   OUT   std_logic;
      DO20                        :   OUT   std_logic;
      DO21                        :   OUT   std_logic;
      DO22                        :   OUT   std_logic;
      DO23                        :   OUT   std_logic;
      DO24                        :   OUT   std_logic;
      DO25                        :   OUT   std_logic;
      DO26                        :   OUT   std_logic;
      DO27                        :   OUT   std_logic;
      DO28                        :   OUT   std_logic;
      DO29                        :   OUT   std_logic;
      DO30                        :   OUT   std_logic;
      DO31                        :   OUT   std_logic;
      DO32                        :   OUT   std_logic;
      DO33                        :   OUT   std_logic;
      DO34                        :   OUT   std_logic;
      DO35                        :   OUT   std_logic;
      DO36                        :   OUT   std_logic;
      DO37                        :   OUT   std_logic;
      DO38                        :   OUT   std_logic;
      DO39                        :   OUT   std_logic;
      DO40                        :   OUT   std_logic;
      DO41                        :   OUT   std_logic;
      DO42                        :   OUT   std_logic;
      DO43                        :   OUT   std_logic;
      DO44                        :   OUT   std_logic;
      DO45                        :   OUT   std_logic;
      DO46                        :   OUT   std_logic;
      DO47                        :   OUT   std_logic;
      DO48                        :   OUT   std_logic;
      DO49                        :   OUT   std_logic;
      DO50                        :   OUT   std_logic;
      DO51                        :   OUT   std_logic;
      DO52                        :   OUT   std_logic;
      DO53                        :   OUT   std_logic;
      DO54                        :   OUT   std_logic;
      DO55                        :   OUT   std_logic;
      DO56                        :   OUT   std_logic;
      DO57                        :   OUT   std_logic;
      DO58                        :   OUT   std_logic;
      DO59                        :   OUT   std_logic;
      DO60                        :   OUT   std_logic;
      DO61                        :   OUT   std_logic;
      DO62                        :   OUT   std_logic;
      DO63                        :   OUT   std_logic;
      DO64                        :   OUT   std_logic;
      DO65                        :   OUT   std_logic;
      DO66                        :   OUT   std_logic;
      DO67                        :   OUT   std_logic;
      DO68                        :   OUT   std_logic;
      DO69                        :   OUT   std_logic;
      DO70                        :   OUT   std_logic;
      DO71                        :   OUT   std_logic;
      DO72                        :   OUT   std_logic;
      DO73                        :   OUT   std_logic;
      DO74                        :   OUT   std_logic;
      DO75                        :   OUT   std_logic;
      DO76                        :   OUT   std_logic;
      DO77                        :   OUT   std_logic;
      DO78                        :   OUT   std_logic;
      DO79                        :   OUT   std_logic;
      DO80                        :   OUT   std_logic;
      DO81                        :   OUT   std_logic;
      DO82                        :   OUT   std_logic;
      DO83                        :   OUT   std_logic;
      DO84                        :   OUT   std_logic;
      DO85                        :   OUT   std_logic;
      DO86                        :   OUT   std_logic;
      DO87                        :   OUT   std_logic;
      DO88                        :   OUT   std_logic;
      DO89                        :   OUT   std_logic;
      DO90                        :   OUT   std_logic;
      DO91                        :   OUT   std_logic;
      DO92                        :   OUT   std_logic;
      DO93                        :   OUT   std_logic;
      DO94                        :   OUT   std_logic;
      DO95                        :   OUT   std_logic;
      DO96                        :   OUT   std_logic;
      DO97                        :   OUT   std_logic;
      DO98                        :   OUT   std_logic;
      DO99                        :   OUT   std_logic;
      DO100                       :   OUT   std_logic;
      DO101                       :   OUT   std_logic;
      DO102                       :   OUT   std_logic;
      DO103                       :   OUT   std_logic;
      DO104                       :   OUT   std_logic;
      DO105                       :   OUT   std_logic;
      DO106                       :   OUT   std_logic;
      DO107                       :   OUT   std_logic;
      DO108                       :   OUT   std_logic;
      DO109                       :   OUT   std_logic;
      DO110                       :   OUT   std_logic;
      DO111                       :   OUT   std_logic;
      DO112                       :   OUT   std_logic;
      DO113                       :   OUT   std_logic;
      DO114                       :   OUT   std_logic;
      DO115                       :   OUT   std_logic;
      DO116                       :   OUT   std_logic;
      DO117                       :   OUT   std_logic;
      DO118                       :   OUT   std_logic;
      DO119                       :   OUT   std_logic;
      DO120                       :   OUT   std_logic;
      DO121                       :   OUT   std_logic;
      DO122                       :   OUT   std_logic;
      DO123                       :   OUT   std_logic;
      DO124                       :   OUT   std_logic;
      DO125                       :   OUT   std_logic;
      DO126                       :   OUT   std_logic;
      DO127                       :   OUT   std_logic;
      DI0                         :   IN   std_logic;
      DI1                         :   IN   std_logic;
      DI2                         :   IN   std_logic;
      DI3                         :   IN   std_logic;
      DI4                         :   IN   std_logic;
      DI5                         :   IN   std_logic;
      DI6                         :   IN   std_logic;
      DI7                         :   IN   std_logic;
      DI8                         :   IN   std_logic;
      DI9                         :   IN   std_logic;
      DI10                        :   IN   std_logic;
      DI11                        :   IN   std_logic;
      DI12                        :   IN   std_logic;
      DI13                        :   IN   std_logic;
      DI14                        :   IN   std_logic;
      DI15                        :   IN   std_logic;
      DI16                        :   IN   std_logic;
      DI17                        :   IN   std_logic;
      DI18                        :   IN   std_logic;
      DI19                        :   IN   std_logic;
      DI20                        :   IN   std_logic;
      DI21                        :   IN   std_logic;
      DI22                        :   IN   std_logic;
      DI23                        :   IN   std_logic;
      DI24                        :   IN   std_logic;
      DI25                        :   IN   std_logic;
      DI26                        :   IN   std_logic;
      DI27                        :   IN   std_logic;
      DI28                        :   IN   std_logic;
      DI29                        :   IN   std_logic;
      DI30                        :   IN   std_logic;
      DI31                        :   IN   std_logic;
      DI32                        :   IN   std_logic;
      DI33                        :   IN   std_logic;
      DI34                        :   IN   std_logic;
      DI35                        :   IN   std_logic;
      DI36                        :   IN   std_logic;
      DI37                        :   IN   std_logic;
      DI38                        :   IN   std_logic;
      DI39                        :   IN   std_logic;
      DI40                        :   IN   std_logic;
      DI41                        :   IN   std_logic;
      DI42                        :   IN   std_logic;
      DI43                        :   IN   std_logic;
      DI44                        :   IN   std_logic;
      DI45                        :   IN   std_logic;
      DI46                        :   IN   std_logic;
      DI47                        :   IN   std_logic;
      DI48                        :   IN   std_logic;
      DI49                        :   IN   std_logic;
      DI50                        :   IN   std_logic;
      DI51                        :   IN   std_logic;
      DI52                        :   IN   std_logic;
      DI53                        :   IN   std_logic;
      DI54                        :   IN   std_logic;
      DI55                        :   IN   std_logic;
      DI56                        :   IN   std_logic;
      DI57                        :   IN   std_logic;
      DI58                        :   IN   std_logic;
      DI59                        :   IN   std_logic;
      DI60                        :   IN   std_logic;
      DI61                        :   IN   std_logic;
      DI62                        :   IN   std_logic;
      DI63                        :   IN   std_logic;
      DI64                        :   IN   std_logic;
      DI65                        :   IN   std_logic;
      DI66                        :   IN   std_logic;
      DI67                        :   IN   std_logic;
      DI68                        :   IN   std_logic;
      DI69                        :   IN   std_logic;
      DI70                        :   IN   std_logic;
      DI71                        :   IN   std_logic;
      DI72                        :   IN   std_logic;
      DI73                        :   IN   std_logic;
      DI74                        :   IN   std_logic;
      DI75                        :   IN   std_logic;
      DI76                        :   IN   std_logic;
      DI77                        :   IN   std_logic;
      DI78                        :   IN   std_logic;
      DI79                        :   IN   std_logic;
      DI80                        :   IN   std_logic;
      DI81                        :   IN   std_logic;
      DI82                        :   IN   std_logic;
      DI83                        :   IN   std_logic;
      DI84                        :   IN   std_logic;
      DI85                        :   IN   std_logic;
      DI86                        :   IN   std_logic;
      DI87                        :   IN   std_logic;
      DI88                        :   IN   std_logic;
      DI89                        :   IN   std_logic;
      DI90                        :   IN   std_logic;
      DI91                        :   IN   std_logic;
      DI92                        :   IN   std_logic;
      DI93                        :   IN   std_logic;
      DI94                        :   IN   std_logic;
      DI95                        :   IN   std_logic;
      DI96                        :   IN   std_logic;
      DI97                        :   IN   std_logic;
      DI98                        :   IN   std_logic;
      DI99                        :   IN   std_logic;
      DI100                       :   IN   std_logic;
      DI101                       :   IN   std_logic;
      DI102                       :   IN   std_logic;
      DI103                       :   IN   std_logic;
      DI104                       :   IN   std_logic;
      DI105                       :   IN   std_logic;
      DI106                       :   IN   std_logic;
      DI107                       :   IN   std_logic;
      DI108                       :   IN   std_logic;
      DI109                       :   IN   std_logic;
      DI110                       :   IN   std_logic;
      DI111                       :   IN   std_logic;
      DI112                       :   IN   std_logic;
      DI113                       :   IN   std_logic;
      DI114                       :   IN   std_logic;
      DI115                       :   IN   std_logic;
      DI116                       :   IN   std_logic;
      DI117                       :   IN   std_logic;
      DI118                       :   IN   std_logic;
      DI119                       :   IN   std_logic;
      DI120                       :   IN   std_logic;
      DI121                       :   IN   std_logic;
      DI122                       :   IN   std_logic;
      DI123                       :   IN   std_logic;
      DI124                       :   IN   std_logic;
      DI125                       :   IN   std_logic;
      DI126                       :   IN   std_logic;
      DI127                       :   IN   std_logic;
      WEB                         :   IN   std_logic;
      CK                          :   IN   std_logic;
      CS                          :   IN   std_logic;
      OE                          :   IN   std_logic
      );
  END component;



  -----------------------------------------------------------------------------
  -- Internal signals driven by (i.e. "output" from) each block
  -----------------------------------------------------------------------------
  signal msdin_i      : std_logic;
  signal mbypass_i    : std_logic;
  signal mreset_i     : std_logic;


  signal halt_en             : std_logic;   --high active, will go to halt state
  signal nap_en              : std_logic;   --high active, will go to nap state
  signal wakeup_lp           : std_logic;  -- From wakeup_lp input IO
  signal poweron_finish      : std_logic;  --
  signal reset_iso           : std_logic;  -- to isolate the pe1_core reset
  signal reset_core_n        : std_logic;  -- to reset pe1_core, low active
  signal nap_rec             : std_logic;  -- will recover from nap mode

  signal lp_pwr_ok       : std_logic;

  -----------------------------------------------------------------------------
  -- pe1_core/peri driven signals
  -----------------------------------------------------------------------------
  -- Signals to other blocks
  signal ddi_vld_c1    : std_logic; --CJ
  signal ddi_vld_c2    : std_logic; --CJ
  signal fast_d        : std_logic;
  --signals to core2
  signal  c2_core2_en   : std_logic;  -- core2 enable
  signal  c2_rsc_n      : std_logic;
  signal  c2_crb_out    : std_logic_vector(7 downto 0);
  signal  c2_crb_sel    : std_logic_vector(3 downto 0);
  signal  c2_en_wdog    : std_logic;
  signal  c2_pup_clk    : std_logic;
  signal  c2_pup_irq    : std_logic_vector(1 downto 0);
  signal  c2_r_size     : std_logic_vector(1 downto 0);
  signal  c2_c_size     : std_logic_vector(1 downto 0);
  signal  c2_t_ras      : std_logic_vector(2 downto 0);
  signal  c2_t_rcd      : std_logic_vector(1 downto 0);
  signal  c2_t_rp       : std_logic_vector(1 downto 0);
  -- to memories signals
  signal c1_mpram_a    : std_logic_vector(7 downto 0);   --Modified by CJ
  signal c1_mpram_d    : std_logic_vector(127 downto 0);     --Modified by CJ
  signal c1_mpram_ce   : std_logic_vector(1 downto 0);
  --signal c1_mpram_oe   : std_logic_vector(1 downto 0);
  signal c1_mpram_we_n : std_logic;
  signal c1_gmem_a     : std_logic_vector(9 downto 0);
  signal c1_gmem_d     : std_logic_vector(7 downto 0);
  signal c1_gmem_ce_n  : std_logic;
  signal c1_gmem_we_n  : std_logic;
  signal short_cycle   : std_logic;
  -- to PADS
  signal mirqout_o     : std_logic;
  signal mckout1_o     : std_logic;
  signal msdout_o      : std_logic;

  -----------------------------------------------------------------------------
  -- signals between pe1_core and peri
  -----------------------------------------------------------------------------
  -- pe1_core driven
  signal dbus        : std_logic_vector(7 downto 0);
  signal dqm_size    : std_logic_vector(1 downto 0);
  -- Peri driven
  signal irq0        : std_logic;
  signal irq1        : std_logic;
  -----------------------------------------------------------------------------
  -- Memory driven signals
  -----------------------------------------------------------------------------
  -- MPROM0, MPROM1, MPRAM0, MPRAM1
  signal c1_mp_q      : std_logic_vector(127 downto 0);
  signal c2_mp_q      : std_logic_vector(127 downto 0);
  -- GMEM
  signal c1_gmem_q    : std_logic_vector(7 downto 0);
  signal c2_gmem_q    : std_logic_vector(7 downto 0);

-------------------------------------------------------------------------------
---------------dual core related----------------------------------------------------------
-------------------------------------------------------------------------------
  signal c1_req_i    : std_logic;  -- Request signal of core1
  signal c1_req_rd_i : std_logic;  -- signal indicate that core1 is reading out request from CMDR fifo.
  signal c1_d_dqi    : std_logic_vector(159 downto 0); -- Data in from processor --CJ
  signal c1_d_dqo    : std_logic_vector(127 downto 0); -- Data out to processor --CJ
  signal c2_req_i    : std_logic;  --Requset signal of pe1_core 2.
  signal c2_req_rd_i : std_logic;  -- signal indicate that core2 is reading out request from CMDR fifo.
  signal c2_d_dqi    : std_logic_vector(159 downto 0); -- Data in from processor
  signal c2_d_dqo    : std_logic_vector(127 downto 0); -- Data out to processor

  signal c2_mpram_a    : std_logic_vector(7 downto 0); --CJ
  signal c2_mpram_d    : std_logic_vector(127 downto 0); --CJ
  signal c2_mpram_ce   : std_logic_vector(1 downto 0);
  --signal c2_mpram_oe   : std_logic_vector(1 downto 0);
  --signal c2_mpram_we_n : std_logic;
  signal c2_gmem_a     : std_logic_vector(9 downto 0);
  signal c2_gmem_d     : std_logic_vector(7 downto 0);
  signal c2_gmem_ce_n  : std_logic;
  signal c2_gmem_we_n  : std_logic;

  signal mp_RAM0_DO  : std_logic_vector (127 downto 0);
  signal mp_RAM0_DI  : std_logic_vector (127 downto 0);
  signal mp_RAM0_A   : std_logic_vector (7 downto 0);
  signal mp_RAM0_WE  : std_logic;
  signal mp_RAM0_WEB : std_logic;
  signal mp_RAM0_CS  : std_logic;

begin



  mreset_i <= MRESET;
  MIRQOUT <= mirqout_o;
  MCKOUT1 <= mckout1_o;
  mbypass_i <= MBYPASS;
  -- SW debug
  msdin_i <= MSDIN;
  MSDOUT <= msdout_o;


  wakeup_lp <= MWAKEUP_LP;
  lp_pwr_ok <= MLP_PWR_OK;

  ddi_vld_c1 <= C1_DDI_VLD;
  ddi_vld_c2 <= C2_DDI_VLD;
  C1_REQ <= c1_req_i;
  c1_req_rd <= c1_req_rd_i;
  C2_req <= c2_req_i;
  c2_req_rd <= c2_req_rd_i;
  C1_REQ_D <=c1_d_dqi;
  C2_REQ_D <= c2_d_dqi;
  c1_d_dqo <= C1_IN_D;
  c2_d_dqo <= C2_IN_D;


  mp_RAM0_WE <= mp_RAM0_CS and not mp_RAM0_WEB;


 -----------------------------------------------------------------------------
 -----------------------------------------------------------------------------
 -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- Instantiation of memories
  -----------------------------------------------------------------------------

ram0_asic_gen : if USE_ASIC_MEMORIES generate
  mpram00a : SNPS_RF_SP_UHS_256x64
        port map (
          Q        => mp_RAM0_DO(63 downto 0),
          ADR      => mp_RAM0_A,
          D        => mp_RAM0_DI(63 downto 0),
          WE       => mp_RAM0_WE,
          ME       => '1',
          CLK      => hclk,
          TEST1    => '0',
          TEST_RNM => '0',
          RME      => '0',
          RM       => (others => '0'),
          WA       => (others => '0'),
          WPULSE   => (others => '0'),
          LS       => '0',
          BC0      => '0',
          BC1      => '0',
          BC2      => '0');

  mpram00b : SNPS_RF_SP_UHS_256x64
        port map (
          Q        => mp_RAM0_DO(127 downto 64),
          ADR      => mp_RAM0_A,
          D        => mp_RAM0_DI(127 downto 64),
          WE       => mp_RAM0_WE,
          ME       => '1',
          CLK      => hclk,
          TEST1    => '0',
          TEST_RNM => '0',
          RME      => '0',
          RM       => (others => '0'),
          WA       => (others => '0'),
          WPULSE   => (others => '0'),
          LS       => '0',
          BC0      => '0',
          BC1      => '0',
          BC2      => '0');
end generate;

ram0_sim_gen : if not USE_ASIC_MEMORIES generate

  mpram00: FPGA_SU180_256X128X1BM1A
  PORT MAP (
      A0          => mp_RAM0_A(0),
      A1          => mp_RAM0_A(1),
      A2          => mp_RAM0_A(2),
      A3          => mp_RAM0_A(3),
      A4          => mp_RAM0_A(4),
      A5          => mp_RAM0_A(5),
      A6          => mp_RAM0_A(6),
      A7          => mp_RAM0_A(7),
      DO0         => mp_RAM0_DO(0),
      DO1         => mp_RAM0_DO(1),
      DO2         => mp_RAM0_DO(2),
      DO3         => mp_RAM0_DO(3),
      DO4         => mp_RAM0_DO(4),
      DO5         => mp_RAM0_DO(5),
      DO6         => mp_RAM0_DO(6),
      DO7         => mp_RAM0_DO(7),
      DO8         => mp_RAM0_DO(8),
      DO9         => mp_RAM0_DO(9),
      DO10        => mp_RAM0_DO(10),
      DO11        => mp_RAM0_DO(11),
      DO12        => mp_RAM0_DO(12),
      DO13        => mp_RAM0_DO(13),
      DO14        => mp_RAM0_DO(14),
      DO15        => mp_RAM0_DO(15),
      DO16        => mp_RAM0_DO(16),
      DO17        => mp_RAM0_DO(17),
      DO18        => mp_RAM0_DO(18),
      DO19        => mp_RAM0_DO(19),
      DO20        => mp_RAM0_DO(20),
      DO21        => mp_RAM0_DO(21),
      DO22        => mp_RAM0_DO(22),
      DO23        => mp_RAM0_DO(23),
      DO24        => mp_RAM0_DO(24),
      DO25        => mp_RAM0_DO(25),
      DO26        => mp_RAM0_DO(26),
      DO27        => mp_RAM0_DO(27),
      DO28        => mp_RAM0_DO(28),
      DO29        => mp_RAM0_DO(29),
      DO30        => mp_RAM0_DO(30),
      DO31        => mp_RAM0_DO(31),
      DO32        => mp_RAM0_DO(32),
      DO33        => mp_RAM0_DO(33),
      DO34        => mp_RAM0_DO(34),
      DO35        => mp_RAM0_DO(35),
      DO36        => mp_RAM0_DO(36),
      DO37        => mp_RAM0_DO(37),
      DO38        => mp_RAM0_DO(38),
      DO39        => mp_RAM0_DO(39),
      DO40        => mp_RAM0_DO(40),
      DO41        => mp_RAM0_DO(41),
      DO42        => mp_RAM0_DO(42),
      DO43        => mp_RAM0_DO(43),
      DO44        => mp_RAM0_DO(44),
      DO45        => mp_RAM0_DO(45),
      DO46        => mp_RAM0_DO(46),
      DO47        => mp_RAM0_DO(47),
      DO48        => mp_RAM0_DO(48),
      DO49        => mp_RAM0_DO(49),
      DO50        => mp_RAM0_DO(50),
      DO51        => mp_RAM0_DO(51),
      DO52        => mp_RAM0_DO(52),
      DO53        => mp_RAM0_DO(53),
      DO54        => mp_RAM0_DO(54),
      DO55        => mp_RAM0_DO(55),
      DO56        => mp_RAM0_DO(56),
      DO57        => mp_RAM0_DO(57),
      DO58        => mp_RAM0_DO(58),
      DO59        => mp_RAM0_DO(59),
      DO60        => mp_RAM0_DO(60),
      DO61        => mp_RAM0_DO(61),
      DO62        => mp_RAM0_DO(62),
      DO63        => mp_RAM0_DO(63),
      DO64        => mp_RAM0_DO(64),
      DO65        => mp_RAM0_DO(65),
      DO66        => mp_RAM0_DO(66),
      DO67        => mp_RAM0_DO(67),
      DO68        => mp_RAM0_DO(68),
      DO69        => mp_RAM0_DO(69),
      DO70        => mp_RAM0_DO(70),
      DO71        => mp_RAM0_DO(71),
      DO72        => mp_RAM0_DO(72),
      DO73        => mp_RAM0_DO(73),
      DO74        => mp_RAM0_DO(74),
      DO75        => mp_RAM0_DO(75),
      DO76        => mp_RAM0_DO(76),
      DO77        => mp_RAM0_DO(77),
      DO78        => mp_RAM0_DO(78),
      DO79        => mp_RAM0_DO(79),
      DO80        => mp_RAM0_DO(80),  --CJ
      DO81        => mp_RAM0_DO(81),  --CJ
      DO82        => mp_RAM0_DO(82),  --CJ
      DO83        => mp_RAM0_DO(83),  --CJ
      DO84        => mp_RAM0_DO(84),  --CJ
      DO85        => mp_RAM0_DO(85),  --CJ
      DO86        => mp_RAM0_DO(86),  --CJ
      DO87        => mp_RAM0_DO(87),  --CJ
      DO88        => mp_RAM0_DO(88),  --CJ
      DO89        => mp_RAM0_DO(89),  --CJ
      DO90        => mp_RAM0_DO(90),  --CJ
      DO91        => mp_RAM0_DO(91),  --CJ
      DO92        => mp_RAM0_DO(92),  --CJ
      DO93        => mp_RAM0_DO(93),  --CJ
      DO94        => mp_RAM0_DO(94),  --CJ
      DO95        => mp_RAM0_DO(95),  --CJ
      DO96        => mp_RAM0_DO(96),  --CJ
      DO97        => mp_RAM0_DO(97),  --CJ
      DO98        => mp_RAM0_DO(98),  --CJ
      DO99        => mp_RAM0_DO(99),  --CJ
      DO100       => mp_RAM0_DO(100), --CJ
      DO101       => mp_RAM0_DO(101), --CJ
      DO102       => mp_RAM0_DO(102), --CJ
      DO103       => mp_RAM0_DO(103), --CJ
      DO104       => mp_RAM0_DO(104), --CJ
      DO105       => mp_RAM0_DO(105), --CJ
      DO106       => mp_RAM0_DO(106), --CJ
      DO107       => mp_RAM0_DO(107), --CJ
      DO108       => mp_RAM0_DO(108), --CJ
      DO109       => mp_RAM0_DO(109), --CJ
      DO110       => mp_RAM0_DO(110), --CJ
      DO111       => mp_RAM0_DO(111), --CJ
      DO112       => mp_RAM0_DO(112), --CJ
      DO113       => mp_RAM0_DO(113), --CJ
      DO114       => mp_RAM0_DO(114), --CJ
      DO115       => mp_RAM0_DO(115), --CJ
      DO116       => mp_RAM0_DO(116), --CJ
      DO117       => mp_RAM0_DO(117), --CJ
      DO118       => mp_RAM0_DO(118), --CJ
      DO119       => mp_RAM0_DO(119), --CJ
      DO120       => mp_RAM0_DO(120), --CJ
      DO121       => mp_RAM0_DO(121), --CJ
      DO122       => mp_RAM0_DO(122), --CJ
      DO123       => mp_RAM0_DO(123), --CJ
      DO124       => mp_RAM0_DO(124), --CJ
      DO125       => mp_RAM0_DO(125), --CJ
      DO126       => mp_RAM0_DO(126), --CJ
      DO127       => mp_RAM0_DO(127), --CJ
      DI0         => mp_RAM0_DI(0),
      DI1         => mp_RAM0_DI(1),
      DI2         => mp_RAM0_DI(2),
      DI3         => mp_RAM0_DI(3),
      DI4         => mp_RAM0_DI(4),
      DI5         => mp_RAM0_DI(5),
      DI6         => mp_RAM0_DI(6),
      DI7         => mp_RAM0_DI(7),
      DI8         => mp_RAM0_DI(8),
      DI9         => mp_RAM0_DI(9),
      DI10        => mp_RAM0_DI(10),
      DI11        => mp_RAM0_DI(11),
      DI12        => mp_RAM0_DI(12),
      DI13        => mp_RAM0_DI(13),
      DI14        => mp_RAM0_DI(14),
      DI15        => mp_RAM0_DI(15),
      DI16        => mp_RAM0_DI(16),
      DI17        => mp_RAM0_DI(17),
      DI18        => mp_RAM0_DI(18),
      DI19        => mp_RAM0_DI(19),
      DI20        => mp_RAM0_DI(20),
      DI21        => mp_RAM0_DI(21),
      DI22        => mp_RAM0_DI(22),
      DI23        => mp_RAM0_DI(23),
      DI24        => mp_RAM0_DI(24),
      DI25        => mp_RAM0_DI(25),
      DI26        => mp_RAM0_DI(26),
      DI27        => mp_RAM0_DI(27),
      DI28        => mp_RAM0_DI(28),
      DI29        => mp_RAM0_DI(29),
      DI30        => mp_RAM0_DI(30),
      DI31        => mp_RAM0_DI(31),
      DI32        => mp_RAM0_DI(32),
      DI33        => mp_RAM0_DI(33),
      DI34        => mp_RAM0_DI(34),
      DI35        => mp_RAM0_DI(35),
      DI36        => mp_RAM0_DI(36),
      DI37        => mp_RAM0_DI(37),
      DI38        => mp_RAM0_DI(38),
      DI39        => mp_RAM0_DI(39),
      DI40        => mp_RAM0_DI(40),
      DI41        => mp_RAM0_DI(41),
      DI42        => mp_RAM0_DI(42),
      DI43        => mp_RAM0_DI(43),
      DI44        => mp_RAM0_DI(44),
      DI45        => mp_RAM0_DI(45),
      DI46        => mp_RAM0_DI(46),
      DI47        => mp_RAM0_DI(47),
      DI48        => mp_RAM0_DI(48),
      DI49        => mp_RAM0_DI(49),
      DI50        => mp_RAM0_DI(50),
      DI51        => mp_RAM0_DI(51),
      DI52        => mp_RAM0_DI(52),
      DI53        => mp_RAM0_DI(53),
      DI54        => mp_RAM0_DI(54),
      DI55        => mp_RAM0_DI(55),
      DI56        => mp_RAM0_DI(56),
      DI57        => mp_RAM0_DI(57),
      DI58        => mp_RAM0_DI(58),
      DI59        => mp_RAM0_DI(59),
      DI60        => mp_RAM0_DI(60),
      DI61        => mp_RAM0_DI(61),
      DI62        => mp_RAM0_DI(62),
      DI63        => mp_RAM0_DI(63),
      DI64        => mp_RAM0_DI(64),
      DI65        => mp_RAM0_DI(65),
      DI66        => mp_RAM0_DI(66),
      DI67        => mp_RAM0_DI(67),
      DI68        => mp_RAM0_DI(68),
      DI69        => mp_RAM0_DI(69),
      DI70        => mp_RAM0_DI(70),
      DI71        => mp_RAM0_DI(71),
      DI72        => mp_RAM0_DI(72),
      DI73        => mp_RAM0_DI(73),
      DI74        => mp_RAM0_DI(74),
      DI75        => mp_RAM0_DI(75),
      DI76        => mp_RAM0_DI(76),
      DI77        => mp_RAM0_DI(77),
      DI78        => mp_RAM0_DI(78),
      DI79        => mp_RAM0_DI(79),
      DI80        => mp_RAM0_DI(80),  --CJ
      DI81        => mp_RAM0_DI(81),  --CJ
      DI82        => mp_RAM0_DI(82),  --CJ
      DI83        => mp_RAM0_DI(83),  --CJ
      DI84        => mp_RAM0_DI(84),  --CJ
      DI85        => mp_RAM0_DI(85),  --CJ
      DI86        => mp_RAM0_DI(86),  --CJ
      DI87        => mp_RAM0_DI(87),  --CJ
      DI88        => mp_RAM0_DI(88),  --CJ
      DI89        => mp_RAM0_DI(89),  --CJ
      DI90        => mp_RAM0_DI(90),  --CJ
      DI91        => mp_RAM0_DI(91),  --CJ
      DI92        => mp_RAM0_DI(92),  --CJ
      DI93        => mp_RAM0_DI(93),  --CJ
      DI94        => mp_RAM0_DI(94),  --CJ
      DI95        => mp_RAM0_DI(95),  --CJ
      DI96        => mp_RAM0_DI(96),  --CJ
      DI97        => mp_RAM0_DI(97),  --CJ
      DI98        => mp_RAM0_DI(98),  --CJ
      DI99        => mp_RAM0_DI(99),  --CJ
      DI100       => mp_RAM0_DI(100), --CJ
      DI101       => mp_RAM0_DI(101), --CJ
      DI102       => mp_RAM0_DI(102), --CJ
      DI103       => mp_RAM0_DI(103), --CJ
      DI104       => mp_RAM0_DI(104), --CJ
      DI105       => mp_RAM0_DI(105), --CJ
      DI106       => mp_RAM0_DI(106), --CJ
      DI107       => mp_RAM0_DI(107), --CJ
      DI108       => mp_RAM0_DI(108), --CJ
      DI109       => mp_RAM0_DI(109), --CJ
      DI110       => mp_RAM0_DI(110), --CJ
      DI111       => mp_RAM0_DI(111), --CJ
      DI112       => mp_RAM0_DI(112), --CJ
      DI113       => mp_RAM0_DI(113), --CJ
      DI114       => mp_RAM0_DI(114), --CJ
      DI115       => mp_RAM0_DI(115), --CJ
      DI116       => mp_RAM0_DI(116), --CJ
      DI117       => mp_RAM0_DI(117), --CJ
      DI118       => mp_RAM0_DI(118), --CJ
      DI119       => mp_RAM0_DI(119), --CJ
      DI120       => mp_RAM0_DI(120), --CJ
      DI121       => mp_RAM0_DI(121), --CJ
      DI122       => mp_RAM0_DI(122), --CJ
      DI123       => mp_RAM0_DI(123), --CJ
      DI124       => mp_RAM0_DI(124), --CJ
      DI125       => mp_RAM0_DI(125), --CJ
      DI126       => mp_RAM0_DI(126), --CJ
      DI127       => mp_RAM0_DI(127), --CJ
      WEB         => mp_RAM0_WEB    ,
      CK          => hclk           ,
      CS          => mp_RAM0_CS     ,
      OE          => std_logic'('1')
      );
end generate;

--  -----------------------------------------------------------------------------
--  -- Real time clock  !!! SEPARATELY POWERED !!!
--  -----------------------------------------------------------------------------
    rtc0: entity work.pe1_rtc
     generic map (
      USE_ASIC_MEMORIES => USE_ASIC_MEMORIES )
     port map(
      pllout         => HCLK          ,
      lp_pwr_ok      => lp_pwr_ok     ,
	    halt_en        => halt_en       ,
      nap_en         => nap_en        ,
      wakeup_lp      => wakeup_lp     ,
      poweron_finish => poweron_finish,
      reset_iso      => reset_iso     ,
      reset_core_n   => reset_core_n  ,
      nap_rec        => nap_rec       ,
      --gmem1
      c1_gmem_a      => c1_gmem_a     ,
      c1_gmem_q      => c1_gmem_q     ,
      c1_gmem_d      => c1_gmem_d     ,
      c1_gmem_we_n   => c1_gmem_we_n  ,
      c1_gmem_ce_n   => c1_gmem_ce_n  ,
      --gmem2
      c2_gmem_a      => c2_gmem_a     ,
      c2_gmem_q      => c2_gmem_q     ,
      c2_gmem_d      => c2_gmem_d     ,
      c2_gmem_we_n   => c2_gmem_we_n  ,
      c2_gmem_ce_n   => c2_gmem_ce_n  ,
      --bmem
      dbus           => dbus          
      );

  -----------------------------------------------------------------------------
  -- pe1_core
  -----------------------------------------------------------------------------
  core1: entity work.pe1_core
    generic map ( USE_ASIC_MEMORIES => USE_ASIC_MEMORIES )
    port map(
    -- Clocks to/from clock block
    clk_p         => HCLK             , --: in  std_logic;  -- PLL clock
    even_c        => even_c           ,
    ready         => C1_RDY           ,
    -- Control outputs to the clock block
    fast_d        => fast_d           , --: out std_logic;  -- clk_d speed select
    -- Power on signal
    pwr_ok        => std_logic'('1')  , --'1',--pwr_ok,  --: in  std_logic;  -- Power is on --change by maning to '1'
	---------------------------------------------------------------------
    -- Memory signals
    ---------------------------------------------------------------------
    -- MPRAM signals
    mpram_a       => c1_mpram_a       , --: out std_logic_vector(13 downto 0);-- Address
    mpram_d       => c1_mpram_d       , --: out std_logic_vector(79 downto 0);-- Data to memory
    mpram_ce      => c1_mpram_ce      , --: out std_logic_vector(1 downto 0); -- Chip enable(active high)
    --mpram_oe      => c1_mpram_oe      , --: out std_logic_vector(1 downto 0); -- Output enable(active high)
    mpram_we_n    => c1_mpram_we_n    , --: out std_logic;                    -- Write enable(active low)
    -- MPROM/MPRAM data out bus
    mp_q          => c1_mp_q          , --: in  std_logic_vector(79 downto 0);-- Data from MPROM/MPRAM
    -- GMEM signals
    gmem_a        => c1_gmem_a        , --: out std_logic_vector(9 downto 0);
    gmem_d        => c1_gmem_d        , --: out std_logic_vector(7 downto 0);
    gmem_q        => c1_gmem_q        , --: in  std_logic_vector(7 downto 0);
    gmem_ce_n     => c1_gmem_ce_n     , --: out std_logic;
    gmem_we_n     => c1_gmem_we_n     , --: out std_logic;

    c2_core2_en   => c2_core2_en      ,
    c2_rsc_n      => c2_rsc_n         ,
    c2_crb_sel    => c2_crb_sel       ,
    c2_crb_out    => c2_crb_out       ,
    c2_en_wdog    => c2_en_wdog       ,
    c2_pup_clk    => c2_pup_clk       ,
    c2_pup_irq    => c2_pup_irq       ,
    c2_r_size     => c2_r_size        ,
    c2_c_size     => c2_c_size        ,
    c2_t_ras      => c2_t_ras         ,
    c2_t_rcd      => c2_t_rcd         ,
    c2_t_rp       => c2_t_rp          ,
    short_cycle   => short_cycle      ,
    exe           => EXE              , --CJ
    resume        => RESUME           , --CJ
    id_number     => c1_ID            , --CJ
    req_c1        => c1_req_i         , --CJ
    req_rd_c1     => c1_req_rd_i      ,
    ack_c1        => C1_ACK           ,
    ddi_vld       => ddi_vld_c1       , --CJ
    -- RTC block signals
    reset_core_n   => reset_core_n    ,
    reset_iso      => reset_iso       ,
    poweron_finish => poweron_finish  ,
    nap_rec        => nap_rec         ,
    halt_en        => halt_en         ,
    nap_en         => nap_en          ,
    --  Signals to/from Peripheral block
    dbus          => dbus             ,--: out std_logic_vector(7 downto 0);
    --pd            => pd_s             ,--: out std_logic_vector(2 downto 0);  -- pl_pd
    --aaddr         => aaddr            ,--: out std_logic_vector(4 downto 0);  -- pl_aaddr
    dqm_size      => dqm_size         ,--: out std_logic_vector(1 downto 0);
    irq0          => irq0             ,--: in  std_logic;  -- Interrupt request 0
    irq1          => irq1             ,--: in  std_logic;  -- Interrupt request 1
    adc_ref2v  	  => open             ,--: out	std_logic;	-- Select 2V internal ADC reference (1V)
---------------------------------------------------------------------
    -- PADS
---------------------------------------------------------------------
    -- Misc. signals
    mreset_i      => mreset_i         , --: in  std_logic;  -- Asynchronous reset input
    mirqout_o     => mirqout_o        , --: out std_logic;  -- Interrupt  request output
    mckout1_o     => mckout1_o        , --: out std_logic;  -- Programmable clock out
    msdin_i       => msdin_i          , --: in  std_logic;  -- Serial data in (debug)
    msdout_o      => msdout_o         , --: out std_logic;  -- Serial data out
    mbypass_i     => mbypass_i        ,--: in  std_logic;  -- bypass PLL
    -- Cluster interface
    din_c         => c1_d_dqo         ,  --: in  std_logic_vector(7 downto 0); -- Data input bus  --in std_logic_vector(127 downto 0);
    dout_c        => c1_d_dqi           --: out std_logic_vector(7 downto 0); -- Data output bus --out std_logic_vector(31 downto 0);
    );
  core2 : entity work.pe1_acore
  generic map ( USE_ASIC_MEMORIES => USE_ASIC_MEMORIES )
  port map(
---------------------------------------------------------------------
    -- Signals to/from other blocks
---------------------------------------------------------------------
    -- Clocks to/from clock block
    clk_p         => HCLK             ,
    even_c        => even_c           ,
    ready         => C2_RDY           ,
    -- signals from the master pe1_core
    rst_cn        => c2_core2_en      ,       --reset core2 if disabled
    rsc_n         => c2_rsc_n         ,
    clkreq_gen    => std_logic'('0')  , --'0',
    id_number     => c2_ID            ,
    core2_en      => c2_core2_en      ,
    crb_out       => c2_crb_out       ,
    en_wdog       => c2_en_wdog       ,
    pup_clk       => c2_pup_clk       ,
    pup_irq    	  => c2_pup_irq    	  ,
    r_size     	  => c2_r_size     	  ,
    c_size     	  => c2_c_size     	  ,
    t_ras      	  => c2_t_ras      	  ,
    t_rcd      	  => c2_t_rcd      	  ,
    t_rp       	  => c2_t_rp       	  ,
    dqm_size      => dqm_size         ,
    fast_d        => fast_d           ,
    short_cycle   => short_cycle      ,

    crb_sel       => c2_crb_sel       ,
    --  Signals to/from Peripheral block
    irq0          => std_logic'('1')  , --'1',  -- Interrupt request 0
    irq1          => std_logic'('1')  , --'1',  -- Interrupt request 1
---------------------------------------------------------------------
    -- Memory signals
---------------------------------------------------------------------
    -- MPRAM signals
    mpram_a       => c2_mpram_a     ,-- Address
    mpram_d       => c2_mpram_d     ,-- Data to memory
    mpram_ce      => c2_mpram_ce    ,-- Chip enable(active high)
    --mpram_oe      => c2_mpram_oe    ,-- Output enable(active high)
    --mpram_we_n    => c2_mpram_we_n  ,-- Write enable(active low)
    -- MPROM/MPRAM data out bus
    mp_q          => c2_mp_q        ,-- Data from MPROM/MPRAM
    -- GMEM signals
    gmem_a        => c2_gmem_a      ,
    gmem_d        => c2_gmem_d      ,
    gmem_q        => c2_gmem_q      ,
    gmem_ce_n     => c2_gmem_ce_n   ,
    gmem_we_n     => c2_gmem_we_n   ,
    exe           => exe            ,     --CJ
    req_c2        => c2_req_i       ,
    req_rd_c2     => c2_req_rd_i    ,
    ack_c2        => C2_ACK         ,
    ddi_vld       =>ddi_vld_c2      , --CJ
    resume        => RESUME         ,   --CJ
    -- Cluster interface
    din_c         => c2_d_dqo   ,   --in std_logic_vector(127 downto 0)-- Data input bus
    dout_c        => c2_d_dqi   -- out std_logic_vector(31 downto 0); -- Data output bus

    );



    mpmem_inf_inst : entity work.pe1_mpmem_inf
  PORT map(
        -- MPRAM signals
        c1_mpram_a     => c1_mpram_a   ,-- Address
        c1_mpram_d     => c1_mpram_d   ,-- Data to memory
        c1_mpram_ce    => c1_mpram_ce  ,-- Chip enable(active high)
        --c1_mpram_oe    => c1_mpram_oe  ,-- Output enable(active high)
        c1_mpram_we_n  => c1_mpram_we_n,-- Write enable(active low)
        c1_mp_q        => c1_mp_q      ,
        -- MPRAM signals
        c2_mpram_a     => c2_mpram_a   ,-- Address
        c2_mpram_d     => c2_mpram_d   ,-- Data to memory
        c2_mpram_ce    => c2_mpram_ce  ,-- Chip enable(active high)
        --c2_mpram_oe    => c2_mpram_oe  ,-- Output enable(active high)
        --c2_mpram_we_n  => c2_mpram_we_n,-- Write enable(active low)
        c2_mp_q        => c2_mp_q      ,
        --RAM0
        RAM0_DO     => mp_RAM0_DO      ,--: in  std_logic_vector (79 downto 0);
        RAM0_DI     => mp_RAM0_DI      ,--: out std_logic_vector (79 downto 0);
        RAM0_A      => mp_RAM0_A       ,--: out std_logic_vector (13 downto 0);
        RAM0_WEB    => mp_RAM0_WEB     ,--: out std_logic;
        RAM0_CS     => mp_RAM0_CS      --: out std_logic;
    );




  -----------------------------------------------------------------------------
  -- Peripherals
  -----------------------------------------------------------------------------
	irq0 <= '1';
	irq1 <= '1';



end struct;