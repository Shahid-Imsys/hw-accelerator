-------------------------------------------------------------------------------
--                                                                           --
--   COPYRIGHT (C)                       Imsys Technologies AB,  2005        --
--                                                                           --
--   The copyright to the document(s) herein is the property of Imsys        --
--   Technologies AB, Sweden.                                                --
--                                                                           --
--   The document(s) may be used and/or copied only with the written         --
--   permission from Imsys Technologies AB or in accordance with the         --
--   terms and conditions stipulated in the agreement/contract under         --
--   which the document(s) have been supplied.                               --
--                                                                           --
-------------------------------------------------------------------------------
-- Title      : req_logic
-- Project    : GP3000
-------------------------------------------------------------------------------
-- File       : Req_logic.vhd
-- Author     : Chuhang Jin
-- Company    : Imsys Technologies AB
-- Date       : 
-------------------------------------------------------------------------------
-- Description: Request buffer logic and data distribution network
--              
--              
-------------------------------------------------------------------------------
-- TO-DO list : 
--              
-------------------------------------------------------------------------------
-- Revisions  :
-- Date                                 Version         Author  Description
-- 2020-10-21                1.0             CJ                 Created
-- 2020-11-15            2.0         CJ         Distribution network added
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.cluster_pkg.all;


entity req_dst_logic is
  generic (USE_ASIC_MEMORIES : boolean := true);
  port(
    --Shared
    CLK_P        : in  std_logic;
    CLK_E        : in  std_logic;       --Generated by PE pair 1 
    EVEN_P       : in  std_logic;
    RESET        : in  std_logic;
    --Requet logic
    REQ_TO_NOC   : out std_logic;
    REQ_SIG      : in  std_logic_vector(15 downto 0);
    REQ_RD_IN    : in  std_logic_vector(15 downto 0);
    ACK_SIG      : out std_logic_vector(15 downto 0);
    PE_REQ_IN    : in  pe_req;          -- pe_req(0) is the last PE (PE 64)
    CMD_OUTPUT   : out std_logic_vector(31 downto 0);   --Command output to CC
    DATA_OUTPUT  : out std_logic_vector(127 downto 0);  --Data output to CC
    RD_FIFO      : in  std_logic;
    FIFO_VLD     : out std_logic;
    --Distribution network
    DATA_VLD     : in  std_logic;
    DATA_NOC     : in  std_logic_vector(127 downto 0);
    PE_UNIT      : in  std_logic_vector(3 downto 0);
    B_CAST       : in  std_logic;
    DATA_VLD_OUT : out std_logic_vector(15 downto 0);
    PE_DATA_OUT  : out pe_data

    );
end entity req_dst_logic;

architecture rtl of req_dst_logic is

  component fifo
    generic(
      DATA_WIDTH         : integer;
      DATA_DEPTH         : integer;
      PROG_FULL_TRESHOLD : integer;
      USE_ASIC_MEMORIES  : boolean := true
      );
    port (
      clk          : in  std_logic;
      --rd_clk : IN STD_LOGIC;
      srst         : in  std_logic;
      din          : in  std_logic_vector(DATA_WIDTH-1 downto 0);
      wr_en        : in  std_logic;
      rd_en        : in  std_logic;
      dout         : out std_logic_vector(DATA_WIDTH-1 downto 0);
      full         : out std_logic;
      almost_full  : out std_logic;
      empty        : out std_logic;
      almost_empty : out std_logic;
      prog_full    : out std_logic;
      valid        : out std_logic;
      counter      : out integer range DATA_DEPTH-1 downto 0
     --wr_rst_busy : OUT STD_LOGIC;
     --rd_rst_busy : OUT STD_LOGIC
      );
  end component;

  signal id_num         : std_logic_vector(3 downto 0)  := "0000";
  signal id_syn         : std_logic_vector(3 downto 0);
  signal id_syn_d       : std_logic_vector(3 downto 0);
  signal poll_act       : std_logic;
  signal fifo_rdy       : std_logic;    --active low
  signal add_in_1       : std_logic_vector(3 downto 0);
  signal add_in_2       : std_logic_vector(3 downto 0)  := "0000";
  signal bs_out         : std_logic_vector(15 downto 0);
  signal pe_mux_out     : std_logic_vector(159 downto 0);
  signal req_core       : std_logic_vector(159 downto 0);
  signal wr             : std_logic;
  signal rd             : std_logic;
  signal full           : std_logic;
  signal almost_full    : std_logic;
  signal empty          : std_logic;
  signal almost_empty   : std_logic;
--    signal wr_req  : std_logic;
  signal ack_sig_i      : std_logic_vector(15 downto 0);  --Will be replaced with a DTM fifo signal.
--    signal loop_c  : integer := 0;
--  signal chain          : std_logic;    --reserved for later use
  signal prog_full_i    : std_logic;
  signal reset_i        : std_logic;
  signal req_to_noc_i   : std_logic;
  signal req_rd_reg     : std_logic_vector(15 downto 0) := (others => '0');
  signal valid_d        : std_logic;
  signal dout_d         : std_logic_vector(159 downto 0);


begin

  reset_i <= not RESET;


-------------------------------------------------------------
--Polling mechanism
-------------------------------------------------------------
--Activation 
  process (clk_p, reset_i)
  begin
    if reset_i = '1' then
      poll_act <= '0';
    elsif rising_edge(clk_p) then
      if fifo_rdy = '0' and req_sig /= (req_sig'range => '0') then
        poll_act <= '1';
        if REQ_RD_IN /= (REQ_RD_IN'range => '0') then
          poll_act <= '0';
        end if;
      else
        poll_act <= '0';
      end if;
    end if;
  end process;


  process(clk_p, reset_i)
  begin
    if reset_i = '1' then
      req_to_noc_i <= '0';
    elsif rising_edge (clk_p) then
      if EVEN_P = '1'then
        if req_rd_reg /= (req_rd_reg'range => '0') then
          req_to_noc_i <= '1';
        else
          req_to_noc_i <= '0';
        end if;
      end if;
    end if;
  end process;
  REQ_TO_NOC <= not empty or req_to_noc_i;
--ID Number Register and write controller
  process(reset_i, poll_act, id_num, req_sig)
  begin
    if reset_i = '1' then
      ack_sig_i <= (others => '0');
    elsif poll_act = '1' then
      ack_sig_i <= (others => '0');     ---handshake ?
      if req_sig(to_integer(15 - unsigned(id_num))) = '1' then
        ack_sig_i(to_integer(unsigned(id_num))) <= '1';
      else
        ack_sig_i(to_integer(unsigned(id_num))) <= '0';
      end if;
    else
      ack_sig_i <= (others => '0');
    end if;
  end process;

  ACK_SIG <= ack_sig_i;

--Barrel Shifter

  process(req_sig, id_num)
    variable sh_0, sh_1, sh_2, sh_3 : std_logic_vector(15 downto 0);
  begin
    sh_3 := req_sig;
    sh_2 := sh_3;
    sh_1 := sh_2;
    sh_0 := sh_1;

    if id_num(3) = '0' then
      sh_3 := req_sig;
    elsif id_num(3) = '1' then
      sh_3 := req_sig(7 downto 0) & req_sig(15 downto 8);
    end if;

    if id_num(2) = '0' then
      sh_2 := sh_3;
    elsif id_num(2) = '1' then
      sh_2 := sh_3(11 downto 0) & sh_3(15 downto 12);
    end if;

    if id_num(1) = '0' then
      sh_1 := sh_2;
    elsif id_num(1) = '1' then
      sh_1 := sh_2(13 downto 0) & sh_2(15 downto 14);
    end if;

    if id_num(0) = '0' then
      sh_0 := sh_1;
    elsif id_num(0) = '1' then
      sh_0 := sh_1(14 downto 0) & sh_1(15);
    end if;

    bs_out <= sh_0;
  end process;

--Priority Encoder 

  process(poll_act, bs_out)
    variable cnt : integer := 0;
  begin
    add_in_2 <= (others => '0');
    if poll_act = '1' then
      cnt := 0;
      for i in 15 downto 0 loop
        if bs_out(i) = '0'then
          cnt := cnt+1;
        elsif bs_out(i) = '1' then
          add_in_2 <= std_logic_vector(to_unsigned(cnt, 4));  --id"0000" is the first PE  
          exit;
        end if;
      end loop;
    end if;
  end process;

--Adder
  add_in_1 <= id_num;
  process(clk_p, reset_i)                        --add_in_2,wr_req,chain,EVEN_P)
  begin
    if reset_i = '1' then
      id_num <= x"0";
    elsif rising_edge(clk_p) then
      if EVEN_P = '1' then              --falling_edge of clk_e, latch id_num
        if REQ_SIG = (REQ_SIG'range => '0') and REQ_RD_IN = (REQ_RD_IN'range => '0') then
          id_num <= x"0";
        else
          if REQ_RD_IN = (REQ_RD_IN'range => '0') then
            id_num <= std_logic_vector(to_unsigned(to_integer(unsigned(add_in_1))+to_integer(unsigned(add_in_2)), 4));
          end if;
        end if;
      end if;
    end if;
  end process;

------synchronize id with request data-------
  process(clk_p, reset_i)
  begin
    if reset_i = '1' then
      id_syn   <= "0000";
      id_syn_d <= "0000";
    elsif rising_edge(clk_p) then
      if EVEN_P = '1' then
        id_syn <= id_num;
      end if;
      id_syn_d <= id_syn;
    end if;
  end process;

----------------------------------------------------------------
--Request Buffer
----------------------------------------------------------------
--PE Mux
  process(clk_p, reset_i)
  begin
    if reset_i = '1' then
      pe_mux_out <= (others => '0');
      req_rd_reg <= (others => '0');
    elsif rising_edge(clk_p) then
      if EVEN_P = '0' then           --rising_edge (clk_e)
        pe_mux_out <= PE_REQ_IN(to_integer(unsigned(id_syn_d)));  --PE req in comes the same clock cycle when req_sig is raised
        req_rd_reg <= REQ_RD_IN;
      end if;
    end if;
  end process;

--Request FIFO
  process(clk_p, reset_i)
  begin
    if reset_i = '1' then
      wr <= '0';
    elsif rising_edge(clk_p)then
      if (req_rd_reg /= (req_rd_reg'range => '0') and EVEN_P = '0') then  --or (wr_req = '1' and EVEN_P = '0')then
        wr <= '1';
      else
        wr <= '0';
      end if;
    end if;
  end process;
--wr <= poll_act;
--Output delay for synchronization with clk_e
  process(clk_p, reset_i)
  begin
    if reset_i = '1' then
      FIFO_VLD    <= '0';
      CMD_OUTPUT  <= (others => '0');
      DATA_OUTPUT <= (others => '0');
    elsif rising_edge(clk_p) then
      FIFO_VLD    <= valid_d;
      CMD_OUTPUT  <= dout_d(159 downto 128);
      DATA_OUTPUT <= dout_d(127 downto 0);
    end if;
  end process;

  req_core <= pe_mux_out;
  fifo_rdy <= almost_full and rd;
  rd       <= RD_FIFO;

----------------------------------------------------------------
--Distribution network
----------------------------------------------------------------
--PE Demux
  process(clk_p, reset_i)  --Should internal destination listed here?
  begin
    if reset_i = '1' then
      DATA_VLD_OUT <= (others => '0');
      pe_data_out  <= (others => (others => '0'));
    elsif rising_edge(clk_p) then
      if EVEN_P = '0' then
        DATA_VLD_OUT <= (others => '0');
        if B_CAST = '1' then
          for i in 15 downto 0 loop
            pe_data_out (i)  <= DATA_NOC;
            DATA_VLD_OUT (i) <= DATA_VLD;
          end loop;
        else
          DATA_VLD_OUT(to_integer(unsigned(PE_UNIT))) <= DATA_VLD;
          pe_data_out(to_integer(unsigned(PE_UNIT)))  <= DATA_NOC;
        end if;
      end if;
    end if;
  end process;

--DATA_VLD_OUT <= data_vld_out_i; 
  request_fifo : fifo
    generic map(
      DATA_WIDTH         => 160,
      DATA_DEPTH         => 1024,
      PROG_FULL_TRESHOLD => 1023,
      USE_ASIC_MEMORIES  => USE_ASIC_MEMORIES
      )
    port map (
      clk          => clk_p,
      --rd_clk => clk_p,
      srst         => reset_i,
      din          => req_core,
      wr_en        => wr,
      rd_en        => rd,
      dout         => dout_d,
      full         => full,
      almost_full  => almost_full,
      empty        => empty,
      almost_empty => almost_empty,
      prog_full    => prog_full_i,
      valid        => valid_d,
      counter      => open
     --wr_rst_busy => open,
     --rd_rst_busy => open
      );

end architecture;
