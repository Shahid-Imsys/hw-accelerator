-- Top entity for Imsys AB Accelerator simulation
-- 
-- Design: Imsys AB
-- Implemented: Bengt Andersson
-- Revision 0


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library work;
use work.defines.all;


entity Accelerator is
	port (
	);
end Accelerator;



architecture struct of Accelerator is


