-- NoC simulation for Imsys Accelerator
-- 
-- Top file
-- Design: Imsys AB
-- Implemented: Bengt Andersson
-- Revision 0

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library work;
use work.defines.all;


entity NoC is
	port (
	);
end NoC;



architecture struct of NoC is

end struct NoC;

