-- GPP simulation for Imsys Accelerator
-- 
-- Top file
-- Design: Imsys AB
-- Implemented: Bengt Andersson
-- Revision 0


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library work;
use work.defines.all;


entity GPP is
	port (
	);
end GPP;



architecture struct of GPP is

end struct GPP;