VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RIIO_EG1D80V_CORNER_45
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CORNER_45 0 0 ;
  SIZE 80 BY 80 ;
  SYMMETRY X Y ;
  SITE corner_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 11.342 53.555 16.402 53.632 ;
        RECT 11.25 53.647 16.356 53.678 ;
        RECT 11.296 53.601 16.356 53.678 ;
        RECT 11.238 53.676 16.31 53.724 ;
        RECT 11.192 53.705 16.264 53.77 ;
        RECT 11.146 53.751 16.218 53.816 ;
        RECT 11.1 53.797 16.172 53.862 ;
        RECT 11.054 53.843 16.126 53.908 ;
        RECT 11.008 53.889 16.08 53.954 ;
        RECT 10.962 53.935 16.034 54 ;
        RECT 10.916 53.981 15.988 54.046 ;
        RECT 10.87 54.027 15.942 54.092 ;
        RECT 10.824 54.073 15.896 54.138 ;
        RECT 10.778 54.119 15.85 54.184 ;
        RECT 10.732 54.165 15.804 54.23 ;
        RECT 10.686 54.211 15.758 54.276 ;
        RECT 10.64 54.257 15.712 54.322 ;
        RECT 10.594 54.303 15.666 54.368 ;
        RECT 10.548 54.349 15.62 54.414 ;
        RECT 10.502 54.395 15.574 54.46 ;
        RECT 10.456 54.441 15.528 54.506 ;
        RECT 10.41 54.487 15.482 54.552 ;
        RECT 10.364 54.533 15.436 54.598 ;
        RECT 10.318 54.579 15.39 54.644 ;
        RECT 10.272 54.625 15.344 54.69 ;
        RECT 10.226 54.671 15.298 54.736 ;
        RECT 10.18 54.717 15.252 54.782 ;
        RECT 10.134 54.763 15.206 54.828 ;
        RECT 10.088 54.809 15.16 54.874 ;
        RECT 10.042 54.855 15.114 54.92 ;
        RECT 9.996 54.901 15.068 54.966 ;
        RECT 9.95 54.947 15.022 55.012 ;
        RECT 9.904 54.993 14.976 55.058 ;
        RECT 9.858 55.039 14.93 55.104 ;
        RECT 9.812 55.085 14.884 55.15 ;
        RECT 9.766 55.131 14.838 55.196 ;
        RECT 9.72 55.177 14.792 55.242 ;
        RECT 9.674 55.223 14.746 55.288 ;
        RECT 9.628 55.269 14.7 55.334 ;
        RECT 9.582 55.315 14.654 55.38 ;
        RECT 9.536 55.361 14.608 55.426 ;
        RECT 9.49 55.407 14.562 55.472 ;
        RECT 9.444 55.453 14.516 55.518 ;
        RECT 9.398 55.499 14.47 55.564 ;
        RECT 9.352 55.545 14.424 55.61 ;
        RECT 9.306 55.591 14.378 55.656 ;
        RECT 9.26 55.637 14.332 55.702 ;
        RECT 9.214 55.683 14.286 55.748 ;
        RECT 9.168 55.729 14.24 55.794 ;
        RECT 9.122 55.775 14.194 55.84 ;
        RECT 9.076 55.821 14.148 55.886 ;
        RECT 9.03 55.867 14.102 55.932 ;
        RECT 8.984 55.913 14.056 55.978 ;
        RECT 8.938 55.959 14.01 56.024 ;
        RECT 8.892 56.005 13.964 56.07 ;
        RECT 8.846 56.051 13.918 56.116 ;
        RECT 8.8 56.097 13.872 56.162 ;
        RECT 8.754 56.143 13.826 56.208 ;
        RECT 8.708 56.189 13.78 56.254 ;
        RECT 8.662 56.235 13.734 56.3 ;
        RECT 8.616 56.281 13.688 56.346 ;
        RECT 8.57 56.327 13.642 56.392 ;
        RECT 8.524 56.373 13.596 56.438 ;
        RECT 8.478 56.419 13.55 56.484 ;
        RECT 8.432 56.465 13.504 56.53 ;
        RECT 8.386 56.511 13.458 56.576 ;
        RECT 8.34 56.557 13.412 56.622 ;
        RECT 8.294 56.603 13.366 56.668 ;
        RECT 8.248 56.649 13.32 56.714 ;
        RECT 8.202 56.695 13.274 56.76 ;
        RECT 8.156 56.741 13.228 56.806 ;
        RECT 8.11 56.787 13.182 56.852 ;
        RECT 8.064 56.833 13.136 56.898 ;
        RECT 8.018 56.879 13.09 56.944 ;
        RECT 7.972 56.925 13.044 56.99 ;
        RECT 7.926 56.971 12.998 57.036 ;
        RECT 7.88 57.017 12.952 57.082 ;
        RECT 7.834 57.063 12.906 57.128 ;
        RECT 7.788 57.109 12.86 57.174 ;
        RECT 7.742 57.155 12.814 57.22 ;
        RECT 7.696 57.201 12.768 57.266 ;
        RECT 7.65 57.247 12.722 57.312 ;
        RECT 7.65 57.247 12.676 57.358 ;
        RECT 7.65 57.247 12.63 57.404 ;
        RECT 7.65 57.247 12.584 57.45 ;
        RECT 7.65 57.247 12.538 57.496 ;
        RECT 7.65 57.247 12.492 57.542 ;
        RECT 7.65 57.247 12.446 57.588 ;
        RECT 7.65 57.247 12.4 57.634 ;
        RECT 7.65 57.247 12.354 57.68 ;
        RECT 7.65 57.247 12.308 57.726 ;
        RECT 7.65 57.247 12.262 57.772 ;
        RECT 7.65 57.247 12.216 57.818 ;
        RECT 7.65 57.247 12.17 57.864 ;
        RECT 7.65 57.247 12.124 57.91 ;
        RECT 7.65 57.247 12.078 57.956 ;
        RECT 7.65 57.247 12.032 58.002 ;
        RECT 7.65 57.247 11.986 58.048 ;
        RECT 7.65 57.247 11.94 58.094 ;
        RECT 7.65 57.247 11.894 58.14 ;
        RECT 7.65 57.247 11.848 58.186 ;
        RECT 7.65 57.247 11.802 58.232 ;
        RECT 7.65 57.247 11.756 58.278 ;
        RECT 7.65 57.247 11.71 58.324 ;
        RECT 7.65 57.247 11.664 58.37 ;
        RECT 7.65 57.247 11.618 58.416 ;
        RECT 7.65 57.247 11.572 58.462 ;
        RECT 7.65 57.247 11.526 58.508 ;
        RECT 7.65 57.247 11.48 58.554 ;
        RECT 7.65 57.247 11.434 58.6 ;
        RECT 7.65 57.247 11.388 58.646 ;
        RECT 7.65 57.247 11.342 58.692 ;
        RECT 7.65 57.247 11.296 58.738 ;
        RECT 7.65 57.247 11.25 80 ;
        RECT 57.27 7.65 80 11.25 ;
        RECT 53.662 11.235 58.761 11.26 ;
        RECT 52.236 12.661 57.316 12.718 ;
        RECT 57.25 7.66 57.27 12.751 ;
        RECT 52.19 12.707 57.25 12.784 ;
        RECT 52.282 12.615 57.362 12.672 ;
        RECT 57.204 7.693 57.25 12.784 ;
        RECT 52.144 12.753 57.204 12.83 ;
        RECT 52.328 12.569 57.408 12.626 ;
        RECT 57.158 7.739 57.204 12.83 ;
        RECT 52.098 12.799 57.158 12.876 ;
        RECT 52.374 12.523 57.454 12.58 ;
        RECT 57.112 7.785 57.158 12.876 ;
        RECT 52.052 12.845 57.112 12.922 ;
        RECT 52.42 12.477 57.5 12.534 ;
        RECT 57.066 7.831 57.112 12.922 ;
        RECT 52.006 12.891 57.066 12.968 ;
        RECT 52.466 12.431 57.546 12.488 ;
        RECT 57.02 7.877 57.066 12.968 ;
        RECT 51.96 12.937 57.02 13.014 ;
        RECT 52.512 12.385 57.592 12.442 ;
        RECT 56.974 7.923 57.02 13.014 ;
        RECT 51.914 12.983 56.974 13.06 ;
        RECT 52.558 12.339 57.638 12.396 ;
        RECT 56.928 7.969 56.974 13.06 ;
        RECT 51.868 13.029 56.928 13.106 ;
        RECT 52.604 12.293 57.684 12.35 ;
        RECT 56.882 8.015 56.928 13.106 ;
        RECT 51.822 13.075 56.882 13.152 ;
        RECT 52.65 12.247 57.73 12.304 ;
        RECT 56.836 8.061 56.882 13.152 ;
        RECT 51.776 13.121 56.836 13.198 ;
        RECT 52.696 12.201 57.776 12.258 ;
        RECT 56.79 8.107 56.836 13.198 ;
        RECT 51.73 13.167 56.79 13.244 ;
        RECT 52.742 12.155 57.822 12.212 ;
        RECT 56.744 8.153 56.79 13.244 ;
        RECT 51.684 13.213 56.744 13.29 ;
        RECT 52.788 12.109 57.868 12.166 ;
        RECT 56.698 8.199 56.744 13.29 ;
        RECT 51.638 13.259 56.698 13.336 ;
        RECT 52.834 12.063 57.914 12.12 ;
        RECT 56.652 8.245 56.698 13.336 ;
        RECT 51.592 13.305 56.652 13.382 ;
        RECT 52.88 12.017 57.96 12.074 ;
        RECT 56.606 8.291 56.652 13.382 ;
        RECT 51.546 13.351 56.606 13.428 ;
        RECT 52.926 11.971 58.006 12.028 ;
        RECT 56.56 8.337 56.606 13.428 ;
        RECT 51.5 13.397 56.56 13.474 ;
        RECT 52.972 11.925 58.052 11.982 ;
        RECT 56.514 8.383 56.56 13.474 ;
        RECT 51.454 13.443 56.514 13.52 ;
        RECT 53.018 11.879 58.098 11.936 ;
        RECT 56.468 8.429 56.514 13.52 ;
        RECT 51.408 13.489 56.468 13.566 ;
        RECT 53.064 11.833 58.144 11.89 ;
        RECT 56.422 8.475 56.468 13.566 ;
        RECT 51.362 13.535 56.422 13.612 ;
        RECT 53.11 11.787 58.19 11.844 ;
        RECT 56.376 8.521 56.422 13.612 ;
        RECT 51.316 13.581 56.376 13.658 ;
        RECT 53.156 11.741 58.236 11.798 ;
        RECT 56.33 8.567 56.376 13.658 ;
        RECT 51.27 13.627 56.33 13.704 ;
        RECT 53.202 11.695 58.282 11.752 ;
        RECT 56.284 8.613 56.33 13.704 ;
        RECT 51.224 13.673 56.284 13.75 ;
        RECT 53.248 11.649 58.328 11.706 ;
        RECT 56.238 8.659 56.284 13.75 ;
        RECT 51.178 13.719 56.238 13.796 ;
        RECT 53.294 11.603 58.374 11.66 ;
        RECT 56.192 8.705 56.238 13.796 ;
        RECT 51.132 13.765 56.192 13.842 ;
        RECT 53.34 11.557 58.42 11.614 ;
        RECT 56.146 8.751 56.192 13.842 ;
        RECT 51.086 13.811 56.146 13.888 ;
        RECT 53.386 11.511 58.466 11.568 ;
        RECT 56.1 8.797 56.146 13.888 ;
        RECT 51.04 13.857 56.1 13.934 ;
        RECT 53.432 11.465 58.512 11.522 ;
        RECT 56.054 8.843 56.1 13.934 ;
        RECT 50.994 13.903 56.054 13.98 ;
        RECT 53.478 11.419 58.558 11.476 ;
        RECT 56.008 8.889 56.054 13.98 ;
        RECT 50.948 13.949 56.008 14.026 ;
        RECT 53.524 11.373 58.604 11.43 ;
        RECT 55.962 8.935 56.008 14.026 ;
        RECT 50.902 13.995 55.962 14.072 ;
        RECT 53.57 11.327 58.65 11.384 ;
        RECT 55.916 8.981 55.962 14.072 ;
        RECT 50.856 14.041 55.916 14.118 ;
        RECT 53.616 11.281 58.696 11.338 ;
        RECT 55.87 9.027 55.916 14.118 ;
        RECT 50.81 14.087 55.87 14.164 ;
        RECT 53.662 11.235 58.742 11.292 ;
        RECT 55.824 9.073 55.87 14.164 ;
        RECT 50.764 14.133 55.824 14.21 ;
        RECT 53.708 11.189 80 11.25 ;
        RECT 55.778 9.119 55.824 14.21 ;
        RECT 50.718 14.179 55.778 14.256 ;
        RECT 53.754 11.143 80 11.25 ;
        RECT 55.732 9.165 55.778 14.256 ;
        RECT 50.672 14.225 55.732 14.302 ;
        RECT 53.8 11.097 80 11.25 ;
        RECT 55.686 9.211 55.732 14.302 ;
        RECT 50.626 14.271 55.686 14.348 ;
        RECT 53.846 11.051 80 11.25 ;
        RECT 55.64 9.257 55.686 14.348 ;
        RECT 50.58 14.317 55.64 14.394 ;
        RECT 53.892 11.005 80 11.25 ;
        RECT 55.594 9.303 55.64 14.394 ;
        RECT 50.534 14.363 55.594 14.44 ;
        RECT 53.938 10.959 80 11.25 ;
        RECT 55.548 9.349 55.594 14.44 ;
        RECT 50.488 14.409 55.548 14.486 ;
        RECT 53.984 10.913 80 11.25 ;
        RECT 55.502 9.395 55.548 14.486 ;
        RECT 50.442 14.455 55.502 14.532 ;
        RECT 54.03 10.867 80 11.25 ;
        RECT 55.456 9.441 55.502 14.532 ;
        RECT 50.396 14.501 55.456 14.578 ;
        RECT 54.076 10.821 80 11.25 ;
        RECT 55.41 9.487 55.456 14.578 ;
        RECT 50.35 14.547 55.41 14.624 ;
        RECT 54.122 10.775 80 11.25 ;
        RECT 55.364 9.533 55.41 14.624 ;
        RECT 50.304 14.593 55.364 14.67 ;
        RECT 54.168 10.729 80 11.25 ;
        RECT 55.318 9.579 55.364 14.67 ;
        RECT 50.258 14.639 55.318 14.716 ;
        RECT 54.214 10.683 80 11.25 ;
        RECT 55.272 9.625 55.318 14.716 ;
        RECT 50.212 14.685 55.272 14.762 ;
        RECT 54.26 10.637 80 11.25 ;
        RECT 55.226 9.671 55.272 14.762 ;
        RECT 50.166 14.731 55.226 14.808 ;
        RECT 54.306 10.591 80 11.25 ;
        RECT 55.18 9.717 55.226 14.808 ;
        RECT 50.12 14.777 55.18 14.854 ;
        RECT 54.352 10.545 80 11.25 ;
        RECT 55.134 9.763 55.18 14.854 ;
        RECT 50.074 14.823 55.134 14.9 ;
        RECT 54.398 10.499 80 11.25 ;
        RECT 55.088 9.809 55.134 14.9 ;
        RECT 50.028 14.869 55.088 14.946 ;
        RECT 54.444 10.453 80 11.25 ;
        RECT 55.042 9.855 55.088 14.946 ;
        RECT 49.982 14.915 55.042 14.992 ;
        RECT 54.49 10.407 80 11.25 ;
        RECT 54.996 9.901 55.042 14.992 ;
        RECT 49.936 14.961 54.996 15.038 ;
        RECT 54.536 10.361 80 11.25 ;
        RECT 54.95 9.947 54.996 15.038 ;
        RECT 49.89 15.007 54.95 15.084 ;
        RECT 54.582 10.315 80 11.25 ;
        RECT 54.904 9.993 54.95 15.084 ;
        RECT 49.844 15.053 54.904 15.13 ;
        RECT 54.628 10.269 80 11.25 ;
        RECT 54.858 10.039 54.904 15.13 ;
        RECT 49.798 15.099 54.858 15.176 ;
        RECT 54.674 10.223 80 11.25 ;
        RECT 54.812 10.085 54.858 15.176 ;
        RECT 49.752 15.145 54.812 15.222 ;
        RECT 54.72 10.177 80 11.25 ;
        RECT 54.766 10.131 54.812 15.222 ;
        RECT 49.706 15.191 54.766 15.268 ;
        RECT 49.66 15.237 54.72 15.314 ;
        RECT 49.614 15.283 54.674 15.36 ;
        RECT 49.568 15.329 54.628 15.406 ;
        RECT 49.522 15.375 54.582 15.452 ;
        RECT 49.476 15.421 54.536 15.498 ;
        RECT 49.43 15.467 54.49 15.544 ;
        RECT 49.384 15.513 54.444 15.59 ;
        RECT 49.338 15.559 54.398 15.636 ;
        RECT 49.292 15.605 54.352 15.682 ;
        RECT 49.246 15.651 54.306 15.728 ;
        RECT 49.2 15.697 54.26 15.774 ;
        RECT 49.154 15.743 54.214 15.82 ;
        RECT 49.108 15.789 54.168 15.866 ;
        RECT 49.062 15.835 54.122 15.912 ;
        RECT 49.016 15.881 54.076 15.958 ;
        RECT 48.97 15.927 54.03 16.004 ;
        RECT 48.924 15.973 53.984 16.05 ;
        RECT 48.878 16.019 53.938 16.096 ;
        RECT 48.832 16.065 53.892 16.142 ;
        RECT 48.786 16.111 53.846 16.188 ;
        RECT 48.74 16.157 53.8 16.234 ;
        RECT 48.694 16.203 53.754 16.28 ;
        RECT 48.648 16.249 53.708 16.326 ;
        RECT 48.602 16.295 53.662 16.372 ;
        RECT 48.556 16.341 53.616 16.418 ;
        RECT 48.51 16.387 53.57 16.464 ;
        RECT 48.464 16.433 53.524 16.51 ;
        RECT 48.418 16.479 53.478 16.556 ;
        RECT 48.372 16.525 53.432 16.602 ;
        RECT 48.326 16.571 53.386 16.648 ;
        RECT 48.28 16.617 53.34 16.694 ;
        RECT 48.234 16.663 53.294 16.74 ;
        RECT 48.188 16.709 53.248 16.786 ;
        RECT 48.142 16.755 53.202 16.832 ;
        RECT 48.096 16.801 53.156 16.878 ;
        RECT 48.05 16.847 53.11 16.924 ;
        RECT 48.004 16.893 53.064 16.97 ;
        RECT 47.958 16.939 53.018 17.016 ;
        RECT 47.912 16.985 52.972 17.062 ;
        RECT 47.866 17.031 52.926 17.108 ;
        RECT 47.82 17.077 52.88 17.154 ;
        RECT 47.774 17.123 52.834 17.2 ;
        RECT 47.728 17.169 52.788 17.246 ;
        RECT 47.682 17.215 52.742 17.292 ;
        RECT 47.636 17.261 52.696 17.338 ;
        RECT 47.59 17.307 52.65 17.384 ;
        RECT 47.544 17.353 52.604 17.43 ;
        RECT 47.498 17.399 52.558 17.476 ;
        RECT 47.452 17.445 52.512 17.522 ;
        RECT 47.406 17.491 52.466 17.568 ;
        RECT 47.36 17.537 52.42 17.614 ;
        RECT 47.314 17.583 52.374 17.66 ;
        RECT 47.268 17.629 52.328 17.706 ;
        RECT 47.222 17.675 52.282 17.752 ;
        RECT 47.176 17.721 52.236 17.798 ;
        RECT 47.13 17.767 52.19 17.844 ;
        RECT 47.084 17.813 52.144 17.89 ;
        RECT 47.038 17.859 52.098 17.936 ;
        RECT 46.992 17.905 52.052 17.982 ;
        RECT 46.946 17.951 52.006 18.028 ;
        RECT 46.9 17.997 51.96 18.074 ;
        RECT 46.854 18.043 51.914 18.12 ;
        RECT 46.808 18.089 51.868 18.166 ;
        RECT 46.762 18.135 51.822 18.212 ;
        RECT 46.716 18.181 51.776 18.258 ;
        RECT 46.67 18.227 51.73 18.304 ;
        RECT 46.624 18.273 51.684 18.35 ;
        RECT 46.578 18.319 51.638 18.396 ;
        RECT 46.532 18.365 51.592 18.442 ;
        RECT 46.486 18.411 51.546 18.488 ;
        RECT 46.44 18.457 51.5 18.534 ;
        RECT 46.394 18.503 51.454 18.58 ;
        RECT 46.348 18.549 51.408 18.626 ;
        RECT 46.302 18.595 51.362 18.672 ;
        RECT 46.256 18.641 51.316 18.718 ;
        RECT 46.21 18.687 51.27 18.764 ;
        RECT 46.164 18.733 51.224 18.81 ;
        RECT 46.118 18.779 51.178 18.856 ;
        RECT 46.072 18.825 51.132 18.902 ;
        RECT 46.026 18.871 51.086 18.948 ;
        RECT 45.98 18.917 51.04 18.994 ;
        RECT 45.934 18.963 50.994 19.04 ;
        RECT 45.888 19.009 50.948 19.086 ;
        RECT 45.842 19.055 50.902 19.132 ;
        RECT 45.796 19.101 50.856 19.178 ;
        RECT 45.75 19.147 50.81 19.224 ;
        RECT 45.704 19.193 50.764 19.27 ;
        RECT 45.658 19.239 50.718 19.316 ;
        RECT 45.612 19.285 50.672 19.362 ;
        RECT 45.566 19.331 50.626 19.408 ;
        RECT 45.52 19.377 50.58 19.454 ;
        RECT 45.474 19.423 50.534 19.5 ;
        RECT 45.428 19.469 50.488 19.546 ;
        RECT 45.382 19.515 50.442 19.592 ;
        RECT 45.336 19.561 50.396 19.638 ;
        RECT 45.29 19.607 50.35 19.684 ;
        RECT 45.244 19.653 50.304 19.73 ;
        RECT 45.198 19.699 50.258 19.776 ;
        RECT 45.152 19.745 50.212 19.822 ;
        RECT 45.106 19.791 50.166 19.868 ;
        RECT 45.06 19.837 50.12 19.914 ;
        RECT 45.014 19.883 50.074 19.96 ;
        RECT 44.968 19.929 50.028 20.006 ;
        RECT 44.922 19.975 49.982 20.052 ;
        RECT 44.876 20.021 49.936 20.098 ;
        RECT 44.83 20.067 49.89 20.144 ;
        RECT 44.784 20.113 49.844 20.19 ;
        RECT 44.738 20.159 49.798 20.236 ;
        RECT 44.692 20.205 49.752 20.282 ;
        RECT 44.646 20.251 49.706 20.328 ;
        RECT 44.6 20.297 49.66 20.374 ;
        RECT 44.554 20.343 49.614 20.42 ;
        RECT 44.508 20.389 49.568 20.466 ;
        RECT 44.462 20.435 49.522 20.512 ;
        RECT 44.416 20.481 49.476 20.558 ;
        RECT 44.37 20.527 49.43 20.604 ;
        RECT 44.324 20.573 49.384 20.65 ;
        RECT 44.278 20.619 49.338 20.696 ;
        RECT 44.232 20.665 49.292 20.742 ;
        RECT 44.186 20.711 49.246 20.788 ;
        RECT 44.14 20.757 49.2 20.834 ;
        RECT 44.094 20.803 49.154 20.88 ;
        RECT 44.048 20.849 49.108 20.926 ;
        RECT 44.002 20.895 49.062 20.972 ;
        RECT 43.956 20.941 49.016 21.018 ;
        RECT 43.91 20.987 48.97 21.064 ;
        RECT 43.864 21.033 48.924 21.11 ;
        RECT 43.818 21.079 48.878 21.156 ;
        RECT 43.772 21.125 48.832 21.202 ;
        RECT 43.726 21.171 48.786 21.248 ;
        RECT 43.68 21.217 48.74 21.294 ;
        RECT 43.634 21.263 48.694 21.34 ;
        RECT 43.588 21.309 48.648 21.386 ;
        RECT 43.542 21.355 48.602 21.432 ;
        RECT 43.496 21.401 48.556 21.478 ;
        RECT 43.45 21.447 48.51 21.524 ;
        RECT 43.404 21.493 48.464 21.57 ;
        RECT 43.358 21.539 48.418 21.616 ;
        RECT 43.312 21.585 48.372 21.662 ;
        RECT 43.266 21.631 48.326 21.708 ;
        RECT 43.22 21.677 48.28 21.754 ;
        RECT 43.174 21.723 48.234 21.8 ;
        RECT 43.128 21.769 48.188 21.846 ;
        RECT 43.082 21.815 48.142 21.892 ;
        RECT 43.036 21.861 48.096 21.938 ;
        RECT 42.99 21.907 48.05 21.984 ;
        RECT 42.944 21.953 48.004 22.03 ;
        RECT 42.898 21.999 47.958 22.076 ;
        RECT 42.852 22.045 47.912 22.122 ;
        RECT 42.806 22.091 47.866 22.168 ;
        RECT 42.76 22.137 47.82 22.214 ;
        RECT 42.714 22.183 47.774 22.26 ;
        RECT 42.668 22.229 47.728 22.306 ;
        RECT 42.622 22.275 47.682 22.352 ;
        RECT 42.576 22.321 47.636 22.398 ;
        RECT 42.53 22.367 47.59 22.444 ;
        RECT 42.484 22.413 47.544 22.49 ;
        RECT 42.438 22.459 47.498 22.536 ;
        RECT 42.392 22.505 47.452 22.582 ;
        RECT 42.346 22.551 47.406 22.628 ;
        RECT 42.3 22.597 47.36 22.674 ;
        RECT 42.254 22.643 47.314 22.72 ;
        RECT 42.208 22.689 47.268 22.766 ;
        RECT 42.162 22.735 47.222 22.812 ;
        RECT 42.116 22.781 47.176 22.858 ;
        RECT 42.07 22.827 47.13 22.904 ;
        RECT 42.024 22.873 47.084 22.95 ;
        RECT 41.978 22.919 47.038 22.996 ;
        RECT 41.932 22.965 46.992 23.042 ;
        RECT 41.886 23.011 46.946 23.088 ;
        RECT 41.84 23.057 46.9 23.134 ;
        RECT 41.794 23.103 46.854 23.18 ;
        RECT 41.748 23.149 46.808 23.226 ;
        RECT 41.702 23.195 46.762 23.272 ;
        RECT 41.656 23.241 46.716 23.318 ;
        RECT 41.61 23.287 46.67 23.364 ;
        RECT 41.564 23.333 46.624 23.41 ;
        RECT 41.518 23.379 46.578 23.456 ;
        RECT 41.472 23.425 46.532 23.502 ;
        RECT 41.426 23.471 46.486 23.548 ;
        RECT 41.38 23.517 46.44 23.594 ;
        RECT 41.334 23.563 46.394 23.64 ;
        RECT 41.288 23.609 46.348 23.686 ;
        RECT 41.242 23.655 46.302 23.732 ;
        RECT 41.196 23.701 46.256 23.778 ;
        RECT 41.15 23.747 46.21 23.824 ;
        RECT 41.104 23.793 46.164 23.87 ;
        RECT 41.058 23.839 46.118 23.916 ;
        RECT 41.012 23.885 46.072 23.962 ;
        RECT 40.966 23.931 46.026 24.008 ;
        RECT 40.92 23.977 45.98 24.054 ;
        RECT 40.874 24.023 45.934 24.1 ;
        RECT 40.828 24.069 45.888 24.146 ;
        RECT 40.782 24.115 45.842 24.192 ;
        RECT 40.736 24.161 45.796 24.238 ;
        RECT 40.69 24.207 45.75 24.284 ;
        RECT 40.644 24.253 45.704 24.33 ;
        RECT 40.598 24.299 45.658 24.376 ;
        RECT 40.552 24.345 45.612 24.422 ;
        RECT 40.506 24.391 45.566 24.468 ;
        RECT 40.46 24.437 45.52 24.514 ;
        RECT 40.414 24.483 45.474 24.56 ;
        RECT 40.368 24.529 45.428 24.606 ;
        RECT 40.322 24.575 45.382 24.652 ;
        RECT 40.276 24.621 45.336 24.698 ;
        RECT 40.23 24.667 45.29 24.744 ;
        RECT 40.184 24.713 45.244 24.79 ;
        RECT 40.138 24.759 45.198 24.836 ;
        RECT 40.092 24.805 45.152 24.882 ;
        RECT 40.046 24.851 45.106 24.928 ;
        RECT 40 24.897 45.06 24.974 ;
        RECT 39.954 24.943 45.014 25.02 ;
        RECT 39.908 24.989 44.968 25.066 ;
        RECT 39.862 25.035 44.922 25.112 ;
        RECT 39.816 25.081 44.876 25.158 ;
        RECT 39.77 25.127 44.83 25.204 ;
        RECT 39.724 25.173 44.784 25.25 ;
        RECT 39.678 25.219 44.738 25.296 ;
        RECT 39.632 25.265 44.692 25.342 ;
        RECT 39.586 25.311 44.646 25.388 ;
        RECT 39.54 25.357 44.6 25.434 ;
        RECT 39.494 25.403 44.554 25.48 ;
        RECT 39.448 25.449 44.508 25.526 ;
        RECT 39.402 25.495 44.462 25.572 ;
        RECT 39.356 25.541 44.416 25.618 ;
        RECT 39.31 25.587 44.37 25.664 ;
        RECT 39.264 25.633 44.324 25.71 ;
        RECT 39.218 25.679 44.278 25.756 ;
        RECT 39.172 25.725 44.232 25.802 ;
        RECT 39.126 25.771 44.186 25.848 ;
        RECT 39.08 25.817 44.14 25.894 ;
        RECT 39.034 25.863 44.094 25.94 ;
        RECT 38.988 25.909 44.048 25.986 ;
        RECT 38.942 25.955 44.002 26.032 ;
        RECT 38.896 26.001 43.956 26.078 ;
        RECT 38.85 26.047 43.91 26.124 ;
        RECT 38.804 26.093 43.864 26.17 ;
        RECT 38.758 26.139 43.818 26.216 ;
        RECT 38.712 26.185 43.772 26.262 ;
        RECT 38.666 26.231 43.726 26.308 ;
        RECT 38.62 26.277 43.68 26.354 ;
        RECT 38.574 26.323 43.634 26.4 ;
        RECT 38.528 26.369 43.588 26.446 ;
        RECT 38.482 26.415 43.542 26.492 ;
        RECT 38.436 26.461 43.496 26.538 ;
        RECT 38.39 26.507 43.45 26.584 ;
        RECT 38.344 26.553 43.404 26.63 ;
        RECT 38.298 26.599 43.358 26.676 ;
        RECT 38.252 26.645 43.312 26.722 ;
        RECT 38.206 26.691 43.266 26.768 ;
        RECT 38.16 26.737 43.22 26.814 ;
        RECT 38.114 26.783 43.174 26.86 ;
        RECT 38.068 26.829 43.128 26.906 ;
        RECT 38.022 26.875 43.082 26.952 ;
        RECT 37.976 26.921 43.036 26.998 ;
        RECT 37.93 26.967 42.99 27.044 ;
        RECT 37.884 27.013 42.944 27.09 ;
        RECT 37.838 27.059 42.898 27.136 ;
        RECT 37.792 27.105 42.852 27.182 ;
        RECT 37.746 27.151 42.806 27.228 ;
        RECT 37.7 27.197 42.76 27.274 ;
        RECT 37.654 27.243 42.714 27.32 ;
        RECT 37.608 27.289 42.668 27.366 ;
        RECT 37.562 27.335 42.622 27.412 ;
        RECT 37.516 27.381 42.576 27.458 ;
        RECT 37.47 27.427 42.53 27.504 ;
        RECT 37.424 27.473 42.484 27.55 ;
        RECT 37.378 27.519 42.438 27.596 ;
        RECT 37.332 27.565 42.392 27.642 ;
        RECT 37.286 27.611 42.346 27.688 ;
        RECT 37.24 27.657 42.3 27.734 ;
        RECT 37.194 27.703 42.254 27.78 ;
        RECT 37.148 27.749 42.208 27.826 ;
        RECT 37.102 27.795 42.162 27.872 ;
        RECT 37.056 27.841 42.116 27.918 ;
        RECT 37.01 27.887 42.07 27.964 ;
        RECT 36.964 27.933 42.024 28.01 ;
        RECT 36.918 27.979 41.978 28.056 ;
        RECT 36.872 28.025 41.932 28.102 ;
        RECT 36.826 28.071 41.886 28.148 ;
        RECT 36.78 28.117 41.84 28.194 ;
        RECT 36.734 28.163 41.794 28.24 ;
        RECT 36.688 28.209 41.748 28.286 ;
        RECT 36.642 28.255 41.702 28.332 ;
        RECT 36.596 28.301 41.656 28.378 ;
        RECT 36.55 28.347 41.61 28.424 ;
        RECT 36.504 28.393 41.564 28.47 ;
        RECT 36.458 28.439 41.518 28.516 ;
        RECT 36.412 28.485 41.472 28.562 ;
        RECT 36.366 28.531 41.426 28.608 ;
        RECT 36.32 28.577 41.38 28.654 ;
        RECT 36.274 28.623 41.334 28.7 ;
        RECT 36.228 28.669 41.288 28.746 ;
        RECT 36.182 28.715 41.242 28.792 ;
        RECT 36.136 28.761 41.196 28.838 ;
        RECT 36.09 28.807 41.15 28.884 ;
        RECT 36.044 28.853 41.104 28.93 ;
        RECT 35.998 28.899 41.058 28.976 ;
        RECT 35.952 28.945 41.012 29.022 ;
        RECT 35.906 28.991 40.966 29.068 ;
        RECT 35.86 29.037 40.92 29.114 ;
        RECT 35.814 29.083 40.874 29.16 ;
        RECT 35.768 29.129 40.828 29.206 ;
        RECT 35.722 29.175 40.782 29.252 ;
        RECT 35.676 29.221 40.736 29.298 ;
        RECT 35.63 29.267 40.69 29.344 ;
        RECT 35.584 29.313 40.644 29.39 ;
        RECT 35.538 29.359 40.598 29.436 ;
        RECT 35.492 29.405 40.552 29.482 ;
        RECT 35.446 29.451 40.506 29.528 ;
        RECT 35.4 29.497 40.46 29.574 ;
        RECT 35.354 29.543 40.414 29.62 ;
        RECT 35.308 29.589 40.368 29.666 ;
        RECT 35.262 29.635 40.322 29.712 ;
        RECT 35.216 29.681 40.276 29.758 ;
        RECT 35.17 29.727 40.23 29.804 ;
        RECT 35.124 29.773 40.184 29.85 ;
        RECT 35.078 29.819 40.138 29.896 ;
        RECT 35.032 29.865 40.092 29.942 ;
        RECT 34.986 29.911 40.046 29.988 ;
        RECT 34.94 29.957 40 30.034 ;
        RECT 34.894 30.003 39.954 30.08 ;
        RECT 34.848 30.049 39.908 30.126 ;
        RECT 34.802 30.095 39.862 30.172 ;
        RECT 34.756 30.141 39.816 30.218 ;
        RECT 34.71 30.187 39.77 30.264 ;
        RECT 34.664 30.233 39.724 30.31 ;
        RECT 34.618 30.279 39.678 30.356 ;
        RECT 34.572 30.325 39.632 30.402 ;
        RECT 34.526 30.371 39.586 30.448 ;
        RECT 34.48 30.417 39.54 30.494 ;
        RECT 34.434 30.463 39.494 30.54 ;
        RECT 34.388 30.509 39.448 30.586 ;
        RECT 34.342 30.555 39.402 30.632 ;
        RECT 34.296 30.601 39.356 30.678 ;
        RECT 34.25 30.647 39.31 30.724 ;
        RECT 34.204 30.693 39.264 30.77 ;
        RECT 34.158 30.739 39.218 30.816 ;
        RECT 34.112 30.785 39.172 30.862 ;
        RECT 34.066 30.831 39.126 30.908 ;
        RECT 34.02 30.877 39.08 30.954 ;
        RECT 33.974 30.923 39.034 31 ;
        RECT 33.928 30.969 38.988 31.046 ;
        RECT 33.882 31.015 38.942 31.092 ;
        RECT 33.836 31.061 38.896 31.138 ;
        RECT 33.79 31.107 38.85 31.184 ;
        RECT 33.744 31.153 38.804 31.23 ;
        RECT 33.698 31.199 38.758 31.276 ;
        RECT 33.652 31.245 38.712 31.322 ;
        RECT 33.606 31.291 38.666 31.368 ;
        RECT 33.56 31.337 38.62 31.414 ;
        RECT 33.514 31.383 38.574 31.46 ;
        RECT 33.468 31.429 38.528 31.506 ;
        RECT 33.422 31.475 38.482 31.552 ;
        RECT 33.376 31.521 38.436 31.598 ;
        RECT 33.33 31.567 38.39 31.644 ;
        RECT 33.284 31.613 38.344 31.69 ;
        RECT 33.238 31.659 38.298 31.736 ;
        RECT 33.192 31.705 38.252 31.782 ;
        RECT 33.146 31.751 38.206 31.828 ;
        RECT 33.1 31.797 38.16 31.874 ;
        RECT 33.054 31.843 38.114 31.92 ;
        RECT 33.008 31.889 38.068 31.966 ;
        RECT 32.962 31.935 38.022 32.012 ;
        RECT 32.916 31.981 37.976 32.058 ;
        RECT 32.87 32.027 37.93 32.104 ;
        RECT 32.824 32.073 37.884 32.15 ;
        RECT 32.778 32.119 37.838 32.196 ;
        RECT 32.732 32.165 37.792 32.242 ;
        RECT 32.686 32.211 37.746 32.288 ;
        RECT 32.64 32.257 37.7 32.334 ;
        RECT 32.594 32.303 37.654 32.38 ;
        RECT 32.548 32.349 37.608 32.426 ;
        RECT 32.502 32.395 37.562 32.472 ;
        RECT 32.456 32.441 37.516 32.518 ;
        RECT 32.41 32.487 37.47 32.564 ;
        RECT 32.364 32.533 37.424 32.61 ;
        RECT 32.318 32.579 37.378 32.656 ;
        RECT 32.272 32.625 37.332 32.702 ;
        RECT 32.226 32.671 37.286 32.748 ;
        RECT 32.18 32.717 37.24 32.794 ;
        RECT 32.134 32.763 37.194 32.84 ;
        RECT 32.088 32.809 37.148 32.886 ;
        RECT 32.042 32.855 37.102 32.932 ;
        RECT 31.996 32.901 37.056 32.978 ;
        RECT 31.95 32.947 37.01 33.024 ;
        RECT 31.904 32.993 36.964 33.07 ;
        RECT 31.858 33.039 36.918 33.116 ;
        RECT 31.812 33.085 36.872 33.162 ;
        RECT 31.766 33.131 36.826 33.208 ;
        RECT 31.72 33.177 36.78 33.254 ;
        RECT 31.674 33.223 36.734 33.3 ;
        RECT 31.628 33.269 36.688 33.346 ;
        RECT 31.582 33.315 36.642 33.392 ;
        RECT 31.536 33.361 36.596 33.438 ;
        RECT 31.49 33.407 36.55 33.484 ;
        RECT 31.444 33.453 36.504 33.53 ;
        RECT 31.398 33.499 36.458 33.576 ;
        RECT 31.352 33.545 36.412 33.622 ;
        RECT 31.306 33.591 36.366 33.668 ;
        RECT 31.26 33.637 36.32 33.714 ;
        RECT 31.214 33.683 36.274 33.76 ;
        RECT 31.168 33.729 36.228 33.806 ;
        RECT 31.122 33.775 36.182 33.852 ;
        RECT 31.076 33.821 36.136 33.898 ;
        RECT 31.03 33.867 36.09 33.944 ;
        RECT 30.984 33.913 36.044 33.99 ;
        RECT 30.938 33.959 35.998 34.036 ;
        RECT 30.892 34.005 35.952 34.082 ;
        RECT 30.846 34.051 35.906 34.128 ;
        RECT 30.8 34.097 35.86 34.174 ;
        RECT 30.754 34.143 35.814 34.22 ;
        RECT 30.708 34.189 35.768 34.266 ;
        RECT 30.662 34.235 35.722 34.312 ;
        RECT 30.616 34.281 35.676 34.358 ;
        RECT 30.57 34.327 35.63 34.404 ;
        RECT 30.524 34.373 35.584 34.45 ;
        RECT 30.478 34.419 35.538 34.496 ;
        RECT 30.432 34.465 35.492 34.542 ;
        RECT 30.386 34.511 35.446 34.588 ;
        RECT 30.34 34.557 35.4 34.634 ;
        RECT 30.294 34.603 35.354 34.68 ;
        RECT 30.248 34.649 35.308 34.726 ;
        RECT 30.202 34.695 35.262 34.772 ;
        RECT 30.156 34.741 35.216 34.818 ;
        RECT 30.11 34.787 35.17 34.864 ;
        RECT 30.064 34.833 35.124 34.91 ;
        RECT 30.018 34.879 35.078 34.956 ;
        RECT 29.972 34.925 35.032 35.002 ;
        RECT 29.926 34.971 34.986 35.048 ;
        RECT 29.88 35.017 34.94 35.094 ;
        RECT 29.834 35.063 34.894 35.14 ;
        RECT 29.788 35.109 34.848 35.186 ;
        RECT 29.742 35.155 34.802 35.232 ;
        RECT 29.696 35.201 34.756 35.278 ;
        RECT 29.65 35.247 34.71 35.324 ;
        RECT 29.604 35.293 34.664 35.37 ;
        RECT 29.558 35.339 34.618 35.416 ;
        RECT 29.512 35.385 34.572 35.462 ;
        RECT 29.466 35.431 34.526 35.508 ;
        RECT 29.42 35.477 34.48 35.554 ;
        RECT 29.374 35.523 34.434 35.6 ;
        RECT 29.328 35.569 34.388 35.646 ;
        RECT 29.282 35.615 34.342 35.692 ;
        RECT 29.236 35.661 34.296 35.738 ;
        RECT 29.19 35.707 34.25 35.784 ;
        RECT 29.144 35.753 34.204 35.83 ;
        RECT 29.098 35.799 34.158 35.876 ;
        RECT 29.052 35.845 34.112 35.922 ;
        RECT 29.006 35.891 34.066 35.968 ;
        RECT 28.96 35.937 34.02 36.014 ;
        RECT 28.914 35.983 33.974 36.06 ;
        RECT 28.868 36.029 33.928 36.106 ;
        RECT 28.822 36.075 33.882 36.152 ;
        RECT 28.776 36.121 33.836 36.198 ;
        RECT 28.73 36.167 33.79 36.244 ;
        RECT 28.684 36.213 33.744 36.29 ;
        RECT 28.638 36.259 33.698 36.336 ;
        RECT 28.592 36.305 33.652 36.382 ;
        RECT 28.546 36.351 33.606 36.428 ;
        RECT 28.5 36.397 33.56 36.474 ;
        RECT 28.454 36.443 33.514 36.52 ;
        RECT 28.408 36.489 33.468 36.566 ;
        RECT 28.362 36.535 33.422 36.612 ;
        RECT 28.316 36.581 33.376 36.658 ;
        RECT 28.27 36.627 33.33 36.704 ;
        RECT 28.224 36.673 33.284 36.75 ;
        RECT 28.178 36.719 33.238 36.796 ;
        RECT 28.132 36.765 33.192 36.842 ;
        RECT 28.086 36.811 33.146 36.888 ;
        RECT 28.04 36.857 33.1 36.934 ;
        RECT 27.994 36.903 33.054 36.98 ;
        RECT 27.948 36.949 33.008 37.026 ;
        RECT 27.902 36.995 32.962 37.072 ;
        RECT 27.856 37.041 32.916 37.118 ;
        RECT 27.81 37.087 32.87 37.164 ;
        RECT 27.764 37.133 32.824 37.21 ;
        RECT 27.718 37.179 32.778 37.256 ;
        RECT 27.672 37.225 32.732 37.302 ;
        RECT 27.626 37.271 32.686 37.348 ;
        RECT 27.58 37.317 32.64 37.394 ;
        RECT 27.534 37.363 32.594 37.44 ;
        RECT 27.488 37.409 32.548 37.486 ;
        RECT 27.442 37.455 32.502 37.532 ;
        RECT 27.396 37.501 32.456 37.578 ;
        RECT 27.35 37.547 32.41 37.624 ;
        RECT 27.304 37.593 32.364 37.67 ;
        RECT 27.258 37.639 32.318 37.716 ;
        RECT 27.212 37.685 32.272 37.762 ;
        RECT 27.166 37.731 32.226 37.808 ;
        RECT 27.12 37.777 32.18 37.854 ;
        RECT 27.074 37.823 32.134 37.9 ;
        RECT 27.028 37.869 32.088 37.946 ;
        RECT 26.982 37.915 32.042 37.992 ;
        RECT 26.936 37.961 31.996 38.038 ;
        RECT 26.89 38.007 31.95 38.084 ;
        RECT 26.844 38.053 31.904 38.13 ;
        RECT 26.798 38.099 31.858 38.176 ;
        RECT 26.752 38.145 31.812 38.222 ;
        RECT 26.706 38.191 31.766 38.268 ;
        RECT 26.66 38.237 31.72 38.314 ;
        RECT 26.614 38.283 31.674 38.36 ;
        RECT 26.568 38.329 31.628 38.406 ;
        RECT 26.522 38.375 31.582 38.452 ;
        RECT 26.476 38.421 31.536 38.498 ;
        RECT 26.43 38.467 31.49 38.544 ;
        RECT 26.384 38.513 31.444 38.59 ;
        RECT 26.338 38.559 31.398 38.636 ;
        RECT 26.292 38.605 31.352 38.682 ;
        RECT 26.246 38.651 31.306 38.728 ;
        RECT 26.2 38.697 31.26 38.774 ;
        RECT 26.154 38.743 31.214 38.82 ;
        RECT 26.108 38.789 31.168 38.866 ;
        RECT 26.062 38.835 31.122 38.912 ;
        RECT 26.016 38.881 31.076 38.958 ;
        RECT 25.97 38.927 31.03 39.004 ;
        RECT 25.924 38.973 30.984 39.05 ;
        RECT 25.878 39.019 30.938 39.096 ;
        RECT 25.832 39.065 30.892 39.142 ;
        RECT 25.786 39.111 30.846 39.188 ;
        RECT 25.74 39.157 30.8 39.234 ;
        RECT 25.694 39.203 30.754 39.28 ;
        RECT 25.648 39.249 30.708 39.326 ;
        RECT 25.602 39.295 30.662 39.372 ;
        RECT 25.556 39.341 30.616 39.418 ;
        RECT 25.51 39.387 30.57 39.464 ;
        RECT 25.464 39.433 30.524 39.51 ;
        RECT 25.418 39.479 30.478 39.556 ;
        RECT 25.372 39.525 30.432 39.602 ;
        RECT 25.326 39.571 30.386 39.648 ;
        RECT 25.28 39.617 30.34 39.694 ;
        RECT 25.234 39.663 30.294 39.74 ;
        RECT 25.188 39.709 30.248 39.786 ;
        RECT 25.142 39.755 30.202 39.832 ;
        RECT 25.096 39.801 30.156 39.878 ;
        RECT 25.05 39.847 30.11 39.924 ;
        RECT 25.004 39.893 30.064 39.97 ;
        RECT 24.958 39.939 30.018 40.016 ;
        RECT 24.912 39.985 29.972 40.062 ;
        RECT 24.866 40.031 29.926 40.108 ;
        RECT 24.82 40.077 29.88 40.154 ;
        RECT 24.774 40.123 29.834 40.2 ;
        RECT 24.728 40.169 29.788 40.246 ;
        RECT 24.682 40.215 29.742 40.292 ;
        RECT 24.636 40.261 29.696 40.338 ;
        RECT 24.59 40.307 29.65 40.384 ;
        RECT 24.544 40.353 29.604 40.43 ;
        RECT 24.498 40.399 29.558 40.476 ;
        RECT 24.452 40.445 29.512 40.522 ;
        RECT 24.406 40.491 29.466 40.568 ;
        RECT 24.36 40.537 29.42 40.614 ;
        RECT 24.314 40.583 29.374 40.66 ;
        RECT 24.268 40.629 29.328 40.706 ;
        RECT 24.222 40.675 29.282 40.752 ;
        RECT 24.176 40.721 29.236 40.798 ;
        RECT 24.13 40.767 29.19 40.844 ;
        RECT 24.084 40.813 29.144 40.89 ;
        RECT 24.038 40.859 29.098 40.936 ;
        RECT 23.992 40.905 29.052 40.982 ;
        RECT 23.946 40.951 29.006 41.028 ;
        RECT 23.9 40.997 28.96 41.074 ;
        RECT 23.854 41.043 28.914 41.12 ;
        RECT 23.808 41.089 28.868 41.166 ;
        RECT 23.762 41.135 28.822 41.212 ;
        RECT 23.716 41.181 28.776 41.258 ;
        RECT 23.67 41.227 28.73 41.304 ;
        RECT 23.624 41.273 28.684 41.35 ;
        RECT 23.578 41.319 28.638 41.396 ;
        RECT 23.532 41.365 28.592 41.442 ;
        RECT 23.486 41.411 28.546 41.488 ;
        RECT 23.44 41.457 28.5 41.534 ;
        RECT 23.394 41.503 28.454 41.58 ;
        RECT 23.348 41.549 28.408 41.626 ;
        RECT 23.302 41.595 28.362 41.672 ;
        RECT 23.256 41.641 28.316 41.718 ;
        RECT 23.21 41.687 28.27 41.764 ;
        RECT 23.164 41.733 28.224 41.81 ;
        RECT 23.118 41.779 28.178 41.856 ;
        RECT 23.072 41.825 28.132 41.902 ;
        RECT 23.026 41.871 28.086 41.948 ;
        RECT 22.98 41.917 28.04 41.994 ;
        RECT 22.934 41.963 27.994 42.04 ;
        RECT 22.888 42.009 27.948 42.086 ;
        RECT 22.842 42.055 27.902 42.132 ;
        RECT 22.796 42.101 27.856 42.178 ;
        RECT 22.75 42.147 27.81 42.224 ;
        RECT 22.704 42.193 27.764 42.27 ;
        RECT 22.658 42.239 27.718 42.316 ;
        RECT 22.612 42.285 27.672 42.362 ;
        RECT 22.566 42.331 27.626 42.408 ;
        RECT 22.52 42.377 27.58 42.454 ;
        RECT 22.474 42.423 27.534 42.5 ;
        RECT 22.428 42.469 27.488 42.546 ;
        RECT 22.382 42.515 27.442 42.592 ;
        RECT 22.336 42.561 27.396 42.638 ;
        RECT 22.29 42.607 27.35 42.684 ;
        RECT 22.244 42.653 27.304 42.73 ;
        RECT 22.198 42.699 27.258 42.776 ;
        RECT 22.152 42.745 27.212 42.822 ;
        RECT 22.106 42.791 27.166 42.868 ;
        RECT 22.06 42.837 27.12 42.914 ;
        RECT 22.014 42.883 27.074 42.96 ;
        RECT 21.968 42.929 27.028 43.006 ;
        RECT 21.922 42.975 26.982 43.052 ;
        RECT 21.876 43.021 26.936 43.098 ;
        RECT 21.83 43.067 26.89 43.144 ;
        RECT 21.784 43.113 26.844 43.19 ;
        RECT 21.738 43.159 26.798 43.236 ;
        RECT 21.692 43.205 26.752 43.282 ;
        RECT 21.646 43.251 26.706 43.328 ;
        RECT 21.6 43.297 26.66 43.374 ;
        RECT 21.554 43.343 26.614 43.42 ;
        RECT 21.508 43.389 26.568 43.466 ;
        RECT 21.462 43.435 26.522 43.512 ;
        RECT 21.416 43.481 26.476 43.558 ;
        RECT 21.37 43.527 26.43 43.604 ;
        RECT 21.324 43.573 26.384 43.65 ;
        RECT 21.278 43.619 26.338 43.696 ;
        RECT 21.232 43.665 26.292 43.742 ;
        RECT 21.186 43.711 26.246 43.788 ;
        RECT 21.14 43.757 26.2 43.834 ;
        RECT 21.094 43.803 26.154 43.88 ;
        RECT 21.048 43.849 26.108 43.926 ;
        RECT 21.002 43.895 26.062 43.972 ;
        RECT 20.956 43.941 26.016 44.018 ;
        RECT 20.91 43.987 25.97 44.064 ;
        RECT 20.864 44.033 25.924 44.11 ;
        RECT 20.818 44.079 25.878 44.156 ;
        RECT 20.772 44.125 25.832 44.202 ;
        RECT 20.726 44.171 25.786 44.248 ;
        RECT 20.68 44.217 25.74 44.294 ;
        RECT 20.634 44.263 25.694 44.34 ;
        RECT 20.588 44.309 25.648 44.386 ;
        RECT 20.542 44.355 25.602 44.432 ;
        RECT 20.496 44.401 25.556 44.478 ;
        RECT 20.45 44.447 25.51 44.524 ;
        RECT 20.404 44.493 25.464 44.57 ;
        RECT 20.358 44.539 25.418 44.616 ;
        RECT 20.312 44.585 25.372 44.662 ;
        RECT 20.266 44.631 25.326 44.708 ;
        RECT 20.22 44.677 25.28 44.754 ;
        RECT 20.174 44.723 25.234 44.8 ;
        RECT 20.128 44.769 25.188 44.846 ;
        RECT 20.082 44.815 25.142 44.892 ;
        RECT 20.036 44.861 25.096 44.938 ;
        RECT 19.99 44.907 25.05 44.984 ;
        RECT 19.944 44.953 25.004 45.03 ;
        RECT 19.898 44.999 24.958 45.076 ;
        RECT 19.852 45.045 24.912 45.122 ;
        RECT 19.806 45.091 24.866 45.168 ;
        RECT 19.76 45.137 24.82 45.214 ;
        RECT 19.714 45.183 24.774 45.26 ;
        RECT 19.668 45.229 24.728 45.306 ;
        RECT 19.622 45.275 24.682 45.352 ;
        RECT 19.576 45.321 24.636 45.398 ;
        RECT 19.53 45.367 24.59 45.444 ;
        RECT 19.484 45.413 24.544 45.49 ;
        RECT 19.438 45.459 24.498 45.536 ;
        RECT 19.392 45.505 24.452 45.582 ;
        RECT 19.346 45.551 24.406 45.628 ;
        RECT 19.3 45.597 24.36 45.674 ;
        RECT 19.254 45.643 24.314 45.72 ;
        RECT 19.208 45.689 24.268 45.766 ;
        RECT 19.162 45.735 24.222 45.812 ;
        RECT 19.116 45.781 24.176 45.858 ;
        RECT 19.07 45.827 24.13 45.904 ;
        RECT 19.024 45.873 24.084 45.95 ;
        RECT 18.978 45.919 24.038 45.996 ;
        RECT 18.932 45.965 23.992 46.042 ;
        RECT 18.886 46.011 23.946 46.088 ;
        RECT 18.84 46.057 23.9 46.134 ;
        RECT 18.794 46.103 23.854 46.18 ;
        RECT 18.748 46.149 23.808 46.226 ;
        RECT 18.702 46.195 23.762 46.272 ;
        RECT 18.656 46.241 23.716 46.318 ;
        RECT 18.61 46.287 23.67 46.364 ;
        RECT 18.564 46.333 23.624 46.41 ;
        RECT 18.518 46.379 23.578 46.456 ;
        RECT 18.472 46.425 23.532 46.502 ;
        RECT 18.426 46.471 23.486 46.548 ;
        RECT 18.38 46.517 23.44 46.594 ;
        RECT 18.334 46.563 23.394 46.64 ;
        RECT 18.288 46.609 23.348 46.686 ;
        RECT 18.242 46.655 23.302 46.732 ;
        RECT 18.196 46.701 23.256 46.778 ;
        RECT 18.15 46.747 23.21 46.824 ;
        RECT 18.104 46.793 23.164 46.87 ;
        RECT 18.058 46.839 23.118 46.916 ;
        RECT 18.012 46.885 23.072 46.962 ;
        RECT 17.966 46.931 23.026 47.008 ;
        RECT 17.92 46.977 22.98 47.054 ;
        RECT 17.874 47.023 22.934 47.1 ;
        RECT 17.828 47.069 22.888 47.146 ;
        RECT 17.782 47.115 22.842 47.192 ;
        RECT 17.736 47.161 22.796 47.238 ;
        RECT 17.69 47.207 22.75 47.284 ;
        RECT 17.644 47.253 22.704 47.33 ;
        RECT 17.598 47.299 22.658 47.376 ;
        RECT 17.552 47.345 22.612 47.422 ;
        RECT 17.506 47.391 22.566 47.468 ;
        RECT 17.46 47.437 22.52 47.514 ;
        RECT 17.414 47.483 22.474 47.56 ;
        RECT 17.368 47.529 22.428 47.606 ;
        RECT 17.322 47.575 22.382 47.652 ;
        RECT 17.276 47.621 22.336 47.698 ;
        RECT 17.23 47.667 22.29 47.744 ;
        RECT 17.184 47.713 22.244 47.79 ;
        RECT 17.138 47.759 22.198 47.836 ;
        RECT 17.092 47.805 22.152 47.882 ;
        RECT 17.046 47.851 22.106 47.928 ;
        RECT 17 47.897 22.06 47.974 ;
        RECT 16.954 47.943 22.014 48.02 ;
        RECT 16.908 47.989 21.968 48.066 ;
        RECT 16.862 48.035 21.922 48.112 ;
        RECT 16.816 48.081 21.876 48.158 ;
        RECT 16.77 48.127 21.83 48.204 ;
        RECT 16.724 48.173 21.784 48.25 ;
        RECT 16.678 48.219 21.738 48.296 ;
        RECT 16.632 48.265 21.692 48.342 ;
        RECT 16.586 48.311 21.646 48.388 ;
        RECT 16.54 48.357 21.6 48.434 ;
        RECT 16.494 48.403 21.554 48.48 ;
        RECT 16.448 48.449 21.508 48.526 ;
        RECT 16.402 48.495 21.462 48.572 ;
        RECT 16.356 48.541 21.416 48.618 ;
        RECT 16.31 48.587 21.37 48.664 ;
        RECT 16.264 48.633 21.324 48.71 ;
        RECT 16.218 48.679 21.278 48.756 ;
        RECT 16.172 48.725 21.232 48.802 ;
        RECT 16.126 48.771 21.186 48.848 ;
        RECT 16.08 48.817 21.14 48.894 ;
        RECT 16.034 48.863 21.094 48.94 ;
        RECT 15.988 48.909 21.048 48.986 ;
        RECT 15.942 48.955 21.002 49.032 ;
        RECT 15.896 49.001 20.956 49.078 ;
        RECT 15.85 49.047 20.91 49.124 ;
        RECT 15.804 49.093 20.864 49.17 ;
        RECT 15.758 49.139 20.818 49.216 ;
        RECT 15.712 49.185 20.772 49.262 ;
        RECT 15.666 49.231 20.726 49.308 ;
        RECT 15.62 49.277 20.68 49.354 ;
        RECT 15.574 49.323 20.634 49.4 ;
        RECT 15.528 49.369 20.588 49.446 ;
        RECT 15.482 49.415 20.542 49.492 ;
        RECT 15.436 49.461 20.496 49.538 ;
        RECT 15.39 49.507 20.45 49.584 ;
        RECT 15.344 49.553 20.404 49.63 ;
        RECT 15.298 49.599 20.358 49.676 ;
        RECT 15.252 49.645 20.312 49.722 ;
        RECT 15.206 49.691 20.266 49.768 ;
        RECT 15.16 49.737 20.22 49.814 ;
        RECT 15.114 49.783 20.174 49.86 ;
        RECT 15.068 49.829 20.128 49.906 ;
        RECT 15.022 49.875 20.082 49.952 ;
        RECT 14.976 49.921 20.036 49.998 ;
        RECT 14.93 49.967 19.99 50.044 ;
        RECT 14.884 50.013 19.944 50.09 ;
        RECT 14.838 50.059 19.898 50.136 ;
        RECT 14.792 50.105 19.852 50.182 ;
        RECT 14.746 50.151 19.806 50.228 ;
        RECT 14.7 50.197 19.76 50.274 ;
        RECT 14.654 50.243 19.714 50.32 ;
        RECT 14.608 50.289 19.668 50.366 ;
        RECT 14.562 50.335 19.622 50.412 ;
        RECT 14.516 50.381 19.576 50.458 ;
        RECT 14.47 50.427 19.53 50.504 ;
        RECT 14.424 50.473 19.484 50.55 ;
        RECT 14.378 50.519 19.438 50.596 ;
        RECT 14.332 50.565 19.392 50.642 ;
        RECT 14.286 50.611 19.346 50.688 ;
        RECT 14.24 50.657 19.3 50.734 ;
        RECT 14.194 50.703 19.254 50.78 ;
        RECT 14.148 50.749 19.208 50.826 ;
        RECT 14.102 50.795 19.162 50.872 ;
        RECT 14.056 50.841 19.116 50.918 ;
        RECT 14.01 50.887 19.07 50.964 ;
        RECT 13.964 50.933 19.024 51.01 ;
        RECT 13.918 50.979 18.978 51.056 ;
        RECT 13.872 51.025 18.932 51.102 ;
        RECT 13.826 51.071 18.886 51.148 ;
        RECT 13.78 51.117 18.84 51.194 ;
        RECT 13.734 51.163 18.794 51.24 ;
        RECT 13.688 51.209 18.748 51.286 ;
        RECT 13.642 51.255 18.702 51.332 ;
        RECT 13.596 51.301 18.656 51.378 ;
        RECT 13.55 51.347 18.61 51.424 ;
        RECT 13.504 51.393 18.564 51.47 ;
        RECT 13.458 51.439 18.518 51.516 ;
        RECT 13.412 51.485 18.472 51.562 ;
        RECT 13.366 51.531 18.426 51.608 ;
        RECT 13.32 51.577 18.38 51.654 ;
        RECT 13.274 51.623 18.334 51.7 ;
        RECT 13.228 51.669 18.288 51.746 ;
        RECT 13.182 51.715 18.242 51.792 ;
        RECT 13.136 51.761 18.196 51.838 ;
        RECT 13.09 51.807 18.15 51.884 ;
        RECT 13.044 51.853 18.104 51.93 ;
        RECT 12.998 51.899 18.058 51.976 ;
        RECT 12.952 51.945 18.012 52.022 ;
        RECT 12.906 51.991 17.966 52.068 ;
        RECT 12.86 52.037 17.92 52.114 ;
        RECT 12.814 52.083 17.874 52.16 ;
        RECT 12.768 52.129 17.828 52.206 ;
        RECT 12.722 52.175 17.782 52.252 ;
        RECT 12.676 52.221 17.736 52.298 ;
        RECT 12.63 52.267 17.69 52.344 ;
        RECT 12.584 52.313 17.644 52.39 ;
        RECT 12.538 52.359 17.598 52.436 ;
        RECT 12.492 52.405 17.552 52.482 ;
        RECT 12.446 52.451 17.506 52.528 ;
        RECT 12.4 52.497 17.46 52.574 ;
        RECT 12.354 52.543 17.414 52.62 ;
        RECT 12.308 52.589 17.368 52.666 ;
        RECT 12.262 52.635 17.322 52.712 ;
        RECT 12.216 52.681 17.276 52.758 ;
        RECT 12.17 52.727 17.23 52.804 ;
        RECT 12.124 52.773 17.184 52.85 ;
        RECT 12.078 52.819 17.138 52.896 ;
        RECT 12.032 52.865 17.092 52.942 ;
        RECT 11.986 52.911 17.046 52.988 ;
        RECT 11.94 52.957 17 53.034 ;
        RECT 11.894 53.003 16.954 53.08 ;
        RECT 11.848 53.049 16.908 53.126 ;
        RECT 11.802 53.095 16.862 53.172 ;
        RECT 11.756 53.141 16.816 53.218 ;
        RECT 11.71 53.187 16.77 53.264 ;
        RECT 11.664 53.233 16.724 53.31 ;
        RECT 11.618 53.279 16.678 53.356 ;
        RECT 11.572 53.325 16.632 53.402 ;
        RECT 11.526 53.371 16.586 53.448 ;
        RECT 11.48 53.417 16.54 53.494 ;
        RECT 11.434 53.463 16.494 53.54 ;
        RECT 11.388 53.509 16.448 53.586 ;
    END
    PORT
      LAYER IB ;
        RECT 56.784 34.705 80 34.75 ;
        RECT 60.362 31.15 80 34.75 ;
        RECT 56.738 34.751 61.853 34.76 ;
        RECT 56.738 34.751 61.834 34.792 ;
        RECT 55.312 36.177 60.362 36.259 ;
        RECT 55.358 36.131 60.408 36.218 ;
        RECT 60.326 31.168 60.362 36.259 ;
        RECT 55.266 36.223 60.326 36.3 ;
        RECT 55.404 36.085 60.454 36.172 ;
        RECT 60.28 31.209 60.326 36.3 ;
        RECT 55.22 36.269 60.28 36.346 ;
        RECT 55.45 36.039 60.5 36.126 ;
        RECT 60.234 31.255 60.28 36.346 ;
        RECT 55.174 36.315 60.234 36.392 ;
        RECT 55.496 35.993 60.546 36.08 ;
        RECT 60.188 31.301 60.234 36.392 ;
        RECT 55.128 36.361 60.188 36.438 ;
        RECT 55.542 35.947 60.592 36.034 ;
        RECT 60.142 31.347 60.188 36.438 ;
        RECT 55.082 36.407 60.142 36.484 ;
        RECT 55.588 35.901 60.638 35.988 ;
        RECT 60.096 31.393 60.142 36.484 ;
        RECT 55.036 36.453 60.096 36.53 ;
        RECT 55.634 35.855 60.684 35.942 ;
        RECT 60.05 31.439 60.096 36.53 ;
        RECT 54.99 36.499 60.05 36.576 ;
        RECT 55.68 35.809 60.73 35.896 ;
        RECT 60.004 31.485 60.05 36.576 ;
        RECT 54.944 36.545 60.004 36.622 ;
        RECT 55.726 35.763 60.776 35.85 ;
        RECT 59.958 31.531 60.004 36.622 ;
        RECT 54.898 36.591 59.958 36.668 ;
        RECT 55.772 35.717 60.822 35.804 ;
        RECT 59.912 31.577 59.958 36.668 ;
        RECT 54.852 36.637 59.912 36.714 ;
        RECT 55.818 35.671 60.868 35.758 ;
        RECT 59.866 31.623 59.912 36.714 ;
        RECT 54.806 36.683 59.866 36.76 ;
        RECT 55.864 35.625 60.914 35.712 ;
        RECT 59.82 31.669 59.866 36.76 ;
        RECT 54.76 36.729 59.82 36.806 ;
        RECT 55.91 35.579 60.96 35.666 ;
        RECT 59.774 31.715 59.82 36.806 ;
        RECT 54.714 36.775 59.774 36.852 ;
        RECT 55.956 35.533 61.006 35.62 ;
        RECT 59.728 31.761 59.774 36.852 ;
        RECT 54.668 36.821 59.728 36.898 ;
        RECT 56.002 35.487 61.052 35.574 ;
        RECT 59.682 31.807 59.728 36.898 ;
        RECT 54.622 36.867 59.682 36.944 ;
        RECT 56.048 35.441 61.098 35.528 ;
        RECT 59.636 31.853 59.682 36.944 ;
        RECT 54.576 36.913 59.636 36.99 ;
        RECT 56.094 35.395 61.144 35.482 ;
        RECT 59.59 31.899 59.636 36.99 ;
        RECT 54.53 36.959 59.59 37.036 ;
        RECT 56.14 35.349 61.19 35.436 ;
        RECT 59.544 31.945 59.59 37.036 ;
        RECT 54.484 37.005 59.544 37.082 ;
        RECT 56.186 35.303 61.236 35.39 ;
        RECT 59.498 31.991 59.544 37.082 ;
        RECT 54.438 37.051 59.498 37.128 ;
        RECT 56.232 35.257 61.282 35.344 ;
        RECT 59.452 32.037 59.498 37.128 ;
        RECT 54.392 37.097 59.452 37.174 ;
        RECT 56.278 35.211 61.328 35.298 ;
        RECT 59.406 32.083 59.452 37.174 ;
        RECT 54.346 37.143 59.406 37.22 ;
        RECT 56.324 35.165 61.374 35.252 ;
        RECT 59.36 32.129 59.406 37.22 ;
        RECT 54.3 37.189 59.36 37.266 ;
        RECT 56.37 35.119 61.42 35.206 ;
        RECT 59.314 32.175 59.36 37.266 ;
        RECT 54.254 37.235 59.314 37.312 ;
        RECT 56.416 35.073 61.466 35.16 ;
        RECT 59.268 32.221 59.314 37.312 ;
        RECT 54.208 37.281 59.268 37.358 ;
        RECT 56.462 35.027 61.512 35.114 ;
        RECT 59.222 32.267 59.268 37.358 ;
        RECT 54.162 37.327 59.222 37.404 ;
        RECT 56.508 34.981 61.558 35.068 ;
        RECT 59.176 32.313 59.222 37.404 ;
        RECT 54.116 37.373 59.176 37.45 ;
        RECT 56.554 34.935 61.604 35.022 ;
        RECT 59.13 32.359 59.176 37.45 ;
        RECT 54.07 37.419 59.13 37.496 ;
        RECT 56.6 34.889 61.65 34.976 ;
        RECT 59.084 32.405 59.13 37.496 ;
        RECT 54.024 37.465 59.084 37.542 ;
        RECT 56.646 34.843 61.696 34.93 ;
        RECT 59.038 32.451 59.084 37.542 ;
        RECT 53.978 37.511 59.038 37.588 ;
        RECT 56.692 34.797 61.742 34.884 ;
        RECT 58.992 32.497 59.038 37.588 ;
        RECT 53.932 37.557 58.992 37.634 ;
        RECT 56.738 34.751 61.788 34.838 ;
        RECT 58.946 32.543 58.992 37.634 ;
        RECT 53.886 37.603 58.946 37.68 ;
        RECT 56.83 34.659 80 34.75 ;
        RECT 58.9 32.589 58.946 37.68 ;
        RECT 53.84 37.649 58.9 37.726 ;
        RECT 56.876 34.613 80 34.75 ;
        RECT 58.854 32.635 58.9 37.726 ;
        RECT 53.794 37.695 58.854 37.772 ;
        RECT 56.922 34.567 80 34.75 ;
        RECT 58.808 32.681 58.854 37.772 ;
        RECT 53.748 37.741 58.808 37.818 ;
        RECT 56.968 34.521 80 34.75 ;
        RECT 58.762 32.727 58.808 37.818 ;
        RECT 53.702 37.787 58.762 37.864 ;
        RECT 57.014 34.475 80 34.75 ;
        RECT 58.716 32.773 58.762 37.864 ;
        RECT 53.656 37.833 58.716 37.91 ;
        RECT 57.06 34.429 80 34.75 ;
        RECT 58.67 32.819 58.716 37.91 ;
        RECT 53.61 37.879 58.67 37.956 ;
        RECT 57.106 34.383 80 34.75 ;
        RECT 58.624 32.865 58.67 37.956 ;
        RECT 53.564 37.925 58.624 38.002 ;
        RECT 57.152 34.337 80 34.75 ;
        RECT 58.578 32.911 58.624 38.002 ;
        RECT 53.518 37.971 58.578 38.048 ;
        RECT 57.198 34.291 80 34.75 ;
        RECT 58.532 32.957 58.578 38.048 ;
        RECT 53.472 38.017 58.532 38.094 ;
        RECT 57.244 34.245 80 34.75 ;
        RECT 58.486 33.003 58.532 38.094 ;
        RECT 53.426 38.063 58.486 38.14 ;
        RECT 57.29 34.199 80 34.75 ;
        RECT 58.44 33.049 58.486 38.14 ;
        RECT 53.38 38.109 58.44 38.186 ;
        RECT 57.336 34.153 80 34.75 ;
        RECT 58.394 33.095 58.44 38.186 ;
        RECT 53.334 38.155 58.394 38.232 ;
        RECT 57.382 34.107 80 34.75 ;
        RECT 58.348 33.141 58.394 38.232 ;
        RECT 53.288 38.201 58.348 38.278 ;
        RECT 57.428 34.061 80 34.75 ;
        RECT 58.302 33.187 58.348 38.278 ;
        RECT 53.242 38.247 58.302 38.324 ;
        RECT 57.474 34.015 80 34.75 ;
        RECT 58.256 33.233 58.302 38.324 ;
        RECT 53.196 38.293 58.256 38.37 ;
        RECT 57.52 33.969 80 34.75 ;
        RECT 58.21 33.279 58.256 38.37 ;
        RECT 53.15 38.339 58.21 38.416 ;
        RECT 57.566 33.923 80 34.75 ;
        RECT 58.164 33.325 58.21 38.416 ;
        RECT 53.104 38.385 58.164 38.462 ;
        RECT 57.612 33.877 80 34.75 ;
        RECT 58.118 33.371 58.164 38.462 ;
        RECT 53.058 38.431 58.118 38.508 ;
        RECT 57.658 33.831 80 34.75 ;
        RECT 58.072 33.417 58.118 38.508 ;
        RECT 53.012 38.477 58.072 38.554 ;
        RECT 57.704 33.785 80 34.75 ;
        RECT 58.026 33.463 58.072 38.554 ;
        RECT 52.966 38.523 58.026 38.6 ;
        RECT 57.75 33.739 80 34.75 ;
        RECT 57.98 33.509 58.026 38.6 ;
        RECT 52.92 38.569 57.98 38.646 ;
        RECT 57.796 33.693 80 34.75 ;
        RECT 57.934 33.555 57.98 38.646 ;
        RECT 52.874 38.615 57.934 38.692 ;
        RECT 57.842 33.647 80 34.75 ;
        RECT 57.888 33.601 57.934 38.692 ;
        RECT 52.828 38.661 57.888 38.738 ;
        RECT 52.782 38.707 57.842 38.784 ;
        RECT 52.736 38.753 57.796 38.83 ;
        RECT 52.69 38.799 57.75 38.876 ;
        RECT 52.644 38.845 57.704 38.922 ;
        RECT 52.598 38.891 57.658 38.968 ;
        RECT 52.552 38.937 57.612 39.014 ;
        RECT 52.506 38.983 57.566 39.06 ;
        RECT 52.46 39.029 57.52 39.106 ;
        RECT 52.414 39.075 57.474 39.152 ;
        RECT 52.368 39.121 57.428 39.198 ;
        RECT 52.322 39.167 57.382 39.244 ;
        RECT 52.276 39.213 57.336 39.29 ;
        RECT 52.23 39.259 57.29 39.336 ;
        RECT 52.184 39.305 57.244 39.382 ;
        RECT 52.138 39.351 57.198 39.428 ;
        RECT 52.092 39.397 57.152 39.474 ;
        RECT 52.046 39.443 57.106 39.52 ;
        RECT 52 39.489 57.06 39.566 ;
        RECT 51.954 39.535 57.014 39.612 ;
        RECT 51.908 39.581 56.968 39.658 ;
        RECT 51.862 39.627 56.922 39.704 ;
        RECT 51.816 39.673 56.876 39.75 ;
        RECT 51.77 39.719 56.83 39.796 ;
        RECT 51.724 39.765 56.784 39.842 ;
        RECT 51.678 39.811 56.738 39.888 ;
        RECT 51.632 39.857 56.692 39.934 ;
        RECT 51.586 39.903 56.646 39.98 ;
        RECT 51.54 39.949 56.6 40.026 ;
        RECT 51.494 39.995 56.554 40.072 ;
        RECT 51.448 40.041 56.508 40.118 ;
        RECT 51.402 40.087 56.462 40.164 ;
        RECT 51.356 40.133 56.416 40.21 ;
        RECT 51.31 40.179 56.37 40.256 ;
        RECT 51.264 40.225 56.324 40.302 ;
        RECT 51.218 40.271 56.278 40.348 ;
        RECT 51.172 40.317 56.232 40.394 ;
        RECT 51.126 40.363 56.186 40.44 ;
        RECT 51.08 40.409 56.14 40.486 ;
        RECT 51.034 40.455 56.094 40.532 ;
        RECT 50.988 40.501 56.048 40.578 ;
        RECT 50.942 40.547 56.002 40.624 ;
        RECT 50.896 40.593 55.956 40.67 ;
        RECT 50.85 40.639 55.91 40.716 ;
        RECT 50.804 40.685 55.864 40.762 ;
        RECT 50.758 40.731 55.818 40.808 ;
        RECT 50.712 40.777 55.772 40.854 ;
        RECT 50.666 40.823 55.726 40.9 ;
        RECT 50.62 40.869 55.68 40.946 ;
        RECT 50.574 40.915 55.634 40.992 ;
        RECT 50.528 40.961 55.588 41.038 ;
        RECT 50.482 41.007 55.542 41.084 ;
        RECT 50.436 41.053 55.496 41.13 ;
        RECT 50.39 41.099 55.45 41.176 ;
        RECT 50.344 41.145 55.404 41.222 ;
        RECT 50.298 41.191 55.358 41.268 ;
        RECT 50.252 41.237 55.312 41.314 ;
        RECT 50.206 41.283 55.266 41.36 ;
        RECT 50.16 41.329 55.22 41.406 ;
        RECT 50.114 41.375 55.174 41.452 ;
        RECT 50.068 41.421 55.128 41.498 ;
        RECT 50.022 41.467 55.082 41.544 ;
        RECT 49.976 41.513 55.036 41.59 ;
        RECT 49.93 41.559 54.99 41.636 ;
        RECT 49.884 41.605 54.944 41.682 ;
        RECT 49.838 41.651 54.898 41.728 ;
        RECT 49.792 41.697 54.852 41.774 ;
        RECT 49.746 41.743 54.806 41.82 ;
        RECT 49.7 41.789 54.76 41.866 ;
        RECT 49.654 41.835 54.714 41.912 ;
        RECT 49.608 41.881 54.668 41.958 ;
        RECT 49.562 41.927 54.622 42.004 ;
        RECT 49.516 41.973 54.576 42.05 ;
        RECT 49.47 42.019 54.53 42.096 ;
        RECT 49.424 42.065 54.484 42.142 ;
        RECT 49.378 42.111 54.438 42.188 ;
        RECT 49.332 42.157 54.392 42.234 ;
        RECT 49.286 42.203 54.346 42.28 ;
        RECT 49.24 42.249 54.3 42.326 ;
        RECT 49.194 42.295 54.254 42.372 ;
        RECT 49.148 42.341 54.208 42.418 ;
        RECT 49.102 42.387 54.162 42.464 ;
        RECT 49.056 42.433 54.116 42.51 ;
        RECT 49.01 42.479 54.07 42.556 ;
        RECT 48.964 42.525 54.024 42.602 ;
        RECT 48.918 42.571 53.978 42.648 ;
        RECT 48.872 42.617 53.932 42.694 ;
        RECT 48.826 42.663 53.886 42.74 ;
        RECT 48.78 42.709 53.84 42.786 ;
        RECT 48.734 42.755 53.794 42.832 ;
        RECT 48.688 42.801 53.748 42.878 ;
        RECT 48.642 42.847 53.702 42.924 ;
        RECT 48.596 42.893 53.656 42.97 ;
        RECT 48.55 42.939 53.61 43.016 ;
        RECT 48.504 42.985 53.564 43.062 ;
        RECT 48.458 43.031 53.518 43.108 ;
        RECT 48.412 43.077 53.472 43.154 ;
        RECT 48.366 43.123 53.426 43.2 ;
        RECT 48.32 43.169 53.38 43.246 ;
        RECT 48.274 43.215 53.334 43.292 ;
        RECT 48.228 43.261 53.288 43.338 ;
        RECT 48.182 43.307 53.242 43.384 ;
        RECT 48.136 43.353 53.196 43.43 ;
        RECT 48.09 43.399 53.15 43.476 ;
        RECT 48.044 43.445 53.104 43.522 ;
        RECT 47.998 43.491 53.058 43.568 ;
        RECT 47.952 43.537 53.012 43.614 ;
        RECT 47.906 43.583 52.966 43.66 ;
        RECT 47.86 43.629 52.92 43.706 ;
        RECT 47.814 43.675 52.874 43.752 ;
        RECT 47.768 43.721 52.828 43.798 ;
        RECT 47.722 43.767 52.782 43.844 ;
        RECT 47.676 43.813 52.736 43.89 ;
        RECT 47.63 43.859 52.69 43.936 ;
        RECT 47.584 43.905 52.644 43.982 ;
        RECT 47.538 43.951 52.598 44.028 ;
        RECT 47.492 43.997 52.552 44.074 ;
        RECT 47.446 44.043 52.506 44.12 ;
        RECT 47.4 44.089 52.46 44.166 ;
        RECT 47.354 44.135 52.414 44.212 ;
        RECT 47.308 44.181 52.368 44.258 ;
        RECT 47.262 44.227 52.322 44.304 ;
        RECT 47.216 44.273 52.276 44.35 ;
        RECT 47.17 44.319 52.23 44.396 ;
        RECT 47.124 44.365 52.184 44.442 ;
        RECT 47.078 44.411 52.138 44.488 ;
        RECT 47.032 44.457 52.092 44.534 ;
        RECT 46.986 44.503 52.046 44.58 ;
        RECT 46.94 44.549 52 44.626 ;
        RECT 46.894 44.595 51.954 44.672 ;
        RECT 46.848 44.641 51.908 44.718 ;
        RECT 46.802 44.687 51.862 44.764 ;
        RECT 46.756 44.733 51.816 44.81 ;
        RECT 46.71 44.779 51.77 44.856 ;
        RECT 46.664 44.825 51.724 44.902 ;
        RECT 46.618 44.871 51.678 44.948 ;
        RECT 46.572 44.917 51.632 44.994 ;
        RECT 46.526 44.963 51.586 45.04 ;
        RECT 46.48 45.009 51.54 45.086 ;
        RECT 46.434 45.055 51.494 45.132 ;
        RECT 46.388 45.101 51.448 45.178 ;
        RECT 46.342 45.147 51.402 45.224 ;
        RECT 46.296 45.193 51.356 45.27 ;
        RECT 46.25 45.239 51.31 45.316 ;
        RECT 46.204 45.285 51.264 45.362 ;
        RECT 46.158 45.331 51.218 45.408 ;
        RECT 46.112 45.377 51.172 45.454 ;
        RECT 46.066 45.423 51.126 45.5 ;
        RECT 46.02 45.469 51.08 45.546 ;
        RECT 45.974 45.515 51.034 45.592 ;
        RECT 45.928 45.561 50.988 45.638 ;
        RECT 45.882 45.607 50.942 45.684 ;
        RECT 45.836 45.653 50.896 45.73 ;
        RECT 45.79 45.699 50.85 45.776 ;
        RECT 45.744 45.745 50.804 45.822 ;
        RECT 45.698 45.791 50.758 45.868 ;
        RECT 45.652 45.837 50.712 45.914 ;
        RECT 45.606 45.883 50.666 45.96 ;
        RECT 45.56 45.929 50.62 46.006 ;
        RECT 45.514 45.975 50.574 46.052 ;
        RECT 45.468 46.021 50.528 46.098 ;
        RECT 45.422 46.067 50.482 46.144 ;
        RECT 45.376 46.113 50.436 46.19 ;
        RECT 45.33 46.159 50.39 46.236 ;
        RECT 45.284 46.205 50.344 46.282 ;
        RECT 45.238 46.251 50.298 46.328 ;
        RECT 45.192 46.297 50.252 46.374 ;
        RECT 45.146 46.343 50.206 46.42 ;
        RECT 45.1 46.389 50.16 46.466 ;
        RECT 45.054 46.435 50.114 46.512 ;
        RECT 45.008 46.481 50.068 46.558 ;
        RECT 44.962 46.527 50.022 46.604 ;
        RECT 44.916 46.573 49.976 46.65 ;
        RECT 44.87 46.619 49.93 46.696 ;
        RECT 44.824 46.665 49.884 46.742 ;
        RECT 44.778 46.711 49.838 46.788 ;
        RECT 44.732 46.757 49.792 46.834 ;
        RECT 44.686 46.803 49.746 46.88 ;
        RECT 44.64 46.849 49.7 46.926 ;
        RECT 44.594 46.895 49.654 46.972 ;
        RECT 44.548 46.941 49.608 47.018 ;
        RECT 44.502 46.987 49.562 47.064 ;
        RECT 44.456 47.033 49.516 47.11 ;
        RECT 44.41 47.079 49.47 47.156 ;
        RECT 44.364 47.125 49.424 47.202 ;
        RECT 44.318 47.171 49.378 47.248 ;
        RECT 44.272 47.217 49.332 47.294 ;
        RECT 44.226 47.263 49.286 47.34 ;
        RECT 44.18 47.309 49.24 47.386 ;
        RECT 44.134 47.355 49.194 47.432 ;
        RECT 44.088 47.401 49.148 47.478 ;
        RECT 44.042 47.447 49.102 47.524 ;
        RECT 43.996 47.493 49.056 47.57 ;
        RECT 43.95 47.539 49.01 47.616 ;
        RECT 43.904 47.585 48.964 47.662 ;
        RECT 43.858 47.631 48.918 47.708 ;
        RECT 43.812 47.677 48.872 47.754 ;
        RECT 43.766 47.723 48.826 47.8 ;
        RECT 43.72 47.769 48.78 47.846 ;
        RECT 43.674 47.815 48.734 47.892 ;
        RECT 43.628 47.861 48.688 47.938 ;
        RECT 43.582 47.907 48.642 47.984 ;
        RECT 43.536 47.953 48.596 48.03 ;
        RECT 43.49 47.999 48.55 48.076 ;
        RECT 43.444 48.045 48.504 48.122 ;
        RECT 43.398 48.091 48.458 48.168 ;
        RECT 43.352 48.137 48.412 48.214 ;
        RECT 43.306 48.183 48.366 48.26 ;
        RECT 43.26 48.229 48.32 48.306 ;
        RECT 43.214 48.275 48.274 48.352 ;
        RECT 43.168 48.321 48.228 48.398 ;
        RECT 43.122 48.367 48.182 48.444 ;
        RECT 43.076 48.413 48.136 48.49 ;
        RECT 43.03 48.459 48.09 48.536 ;
        RECT 42.984 48.505 48.044 48.582 ;
        RECT 42.938 48.551 47.998 48.628 ;
        RECT 42.892 48.597 47.952 48.674 ;
        RECT 42.846 48.643 47.906 48.72 ;
        RECT 42.8 48.689 47.86 48.766 ;
        RECT 42.754 48.735 47.814 48.812 ;
        RECT 42.708 48.781 47.768 48.858 ;
        RECT 42.662 48.827 47.722 48.904 ;
        RECT 42.616 48.873 47.676 48.95 ;
        RECT 42.57 48.919 47.63 48.996 ;
        RECT 42.524 48.965 47.584 49.042 ;
        RECT 42.478 49.011 47.538 49.088 ;
        RECT 42.432 49.057 47.492 49.134 ;
        RECT 42.386 49.103 47.446 49.18 ;
        RECT 42.34 49.149 47.4 49.226 ;
        RECT 42.294 49.195 47.354 49.272 ;
        RECT 42.248 49.241 47.308 49.318 ;
        RECT 42.202 49.287 47.262 49.364 ;
        RECT 42.156 49.333 47.216 49.41 ;
        RECT 42.11 49.379 47.17 49.456 ;
        RECT 42.064 49.425 47.124 49.502 ;
        RECT 42.018 49.471 47.078 49.548 ;
        RECT 41.972 49.517 47.032 49.594 ;
        RECT 41.926 49.563 46.986 49.64 ;
        RECT 41.88 49.609 46.94 49.686 ;
        RECT 41.834 49.655 46.894 49.732 ;
        RECT 41.788 49.701 46.848 49.778 ;
        RECT 41.742 49.747 46.802 49.824 ;
        RECT 41.696 49.793 46.756 49.87 ;
        RECT 41.65 49.839 46.71 49.916 ;
        RECT 41.604 49.885 46.664 49.962 ;
        RECT 41.558 49.931 46.618 50.008 ;
        RECT 41.512 49.977 46.572 50.054 ;
        RECT 41.466 50.023 46.526 50.1 ;
        RECT 41.42 50.069 46.48 50.146 ;
        RECT 41.374 50.115 46.434 50.192 ;
        RECT 41.328 50.161 46.388 50.238 ;
        RECT 41.282 50.207 46.342 50.284 ;
        RECT 41.236 50.253 46.296 50.33 ;
        RECT 41.19 50.299 46.25 50.376 ;
        RECT 41.144 50.345 46.204 50.422 ;
        RECT 41.098 50.391 46.158 50.468 ;
        RECT 41.052 50.437 46.112 50.514 ;
        RECT 41.006 50.483 46.066 50.56 ;
        RECT 40.96 50.529 46.02 50.606 ;
        RECT 40.914 50.575 45.974 50.652 ;
        RECT 40.868 50.621 45.928 50.698 ;
        RECT 40.822 50.667 45.882 50.744 ;
        RECT 40.776 50.713 45.836 50.79 ;
        RECT 40.73 50.759 45.79 50.836 ;
        RECT 40.684 50.805 45.744 50.882 ;
        RECT 40.638 50.851 45.698 50.928 ;
        RECT 40.592 50.897 45.652 50.974 ;
        RECT 40.546 50.943 45.606 51.02 ;
        RECT 40.5 50.989 45.56 51.066 ;
        RECT 40.454 51.035 45.514 51.112 ;
        RECT 40.408 51.081 45.468 51.158 ;
        RECT 40.362 51.127 45.422 51.204 ;
        RECT 40.316 51.173 45.376 51.25 ;
        RECT 40.27 51.219 45.33 51.296 ;
        RECT 40.224 51.265 45.284 51.342 ;
        RECT 40.178 51.311 45.238 51.388 ;
        RECT 40.132 51.357 45.192 51.434 ;
        RECT 40.086 51.403 45.146 51.48 ;
        RECT 40.04 51.449 45.1 51.526 ;
        RECT 39.994 51.495 45.054 51.572 ;
        RECT 39.948 51.541 45.008 51.618 ;
        RECT 39.902 51.587 44.962 51.664 ;
        RECT 39.856 51.633 44.916 51.71 ;
        RECT 39.81 51.679 44.87 51.756 ;
        RECT 39.764 51.725 44.824 51.802 ;
        RECT 39.718 51.771 44.778 51.848 ;
        RECT 39.672 51.817 44.732 51.894 ;
        RECT 39.626 51.863 44.686 51.94 ;
        RECT 39.58 51.909 44.64 51.986 ;
        RECT 39.534 51.955 44.594 52.032 ;
        RECT 39.488 52.001 44.548 52.078 ;
        RECT 39.442 52.047 44.502 52.124 ;
        RECT 39.396 52.093 44.456 52.17 ;
        RECT 39.35 52.139 44.41 52.216 ;
        RECT 39.304 52.185 44.364 52.262 ;
        RECT 39.258 52.231 44.318 52.308 ;
        RECT 39.212 52.277 44.272 52.354 ;
        RECT 39.166 52.323 44.226 52.4 ;
        RECT 39.12 52.369 44.18 52.446 ;
        RECT 39.074 52.415 44.134 52.492 ;
        RECT 39.028 52.461 44.088 52.538 ;
        RECT 38.982 52.507 44.042 52.584 ;
        RECT 38.936 52.553 43.996 52.63 ;
        RECT 38.89 52.599 43.95 52.676 ;
        RECT 38.844 52.645 43.904 52.722 ;
        RECT 38.798 52.691 43.858 52.768 ;
        RECT 38.752 52.737 43.812 52.814 ;
        RECT 38.706 52.783 43.766 52.86 ;
        RECT 38.66 52.829 43.72 52.906 ;
        RECT 38.614 52.875 43.674 52.952 ;
        RECT 38.568 52.921 43.628 52.998 ;
        RECT 38.522 52.967 43.582 53.044 ;
        RECT 38.476 53.013 43.536 53.09 ;
        RECT 38.43 53.059 43.49 53.136 ;
        RECT 38.384 53.105 43.444 53.182 ;
        RECT 38.338 53.151 43.398 53.228 ;
        RECT 38.292 53.197 43.352 53.274 ;
        RECT 38.246 53.243 43.306 53.32 ;
        RECT 38.2 53.289 43.26 53.366 ;
        RECT 38.154 53.335 43.214 53.412 ;
        RECT 38.108 53.381 43.168 53.458 ;
        RECT 38.062 53.427 43.122 53.504 ;
        RECT 38.016 53.473 43.076 53.55 ;
        RECT 37.97 53.519 43.03 53.596 ;
        RECT 37.924 53.565 42.984 53.642 ;
        RECT 37.878 53.611 42.938 53.688 ;
        RECT 37.832 53.657 42.892 53.734 ;
        RECT 37.786 53.703 42.846 53.78 ;
        RECT 37.74 53.749 42.8 53.826 ;
        RECT 37.694 53.795 42.754 53.872 ;
        RECT 37.648 53.841 42.708 53.918 ;
        RECT 37.602 53.887 42.662 53.964 ;
        RECT 37.556 53.933 42.616 54.01 ;
        RECT 37.51 53.979 42.57 54.056 ;
        RECT 37.464 54.025 42.524 54.102 ;
        RECT 37.418 54.071 42.478 54.148 ;
        RECT 37.372 54.117 42.432 54.194 ;
        RECT 37.326 54.163 42.386 54.24 ;
        RECT 37.28 54.209 42.34 54.286 ;
        RECT 37.234 54.255 42.294 54.332 ;
        RECT 37.188 54.301 42.248 54.378 ;
        RECT 37.142 54.347 42.202 54.424 ;
        RECT 37.096 54.393 42.156 54.47 ;
        RECT 37.05 54.439 42.11 54.516 ;
        RECT 37.004 54.485 42.064 54.562 ;
        RECT 36.958 54.531 42.018 54.608 ;
        RECT 36.912 54.577 41.972 54.654 ;
        RECT 36.866 54.623 41.926 54.7 ;
        RECT 36.82 54.669 41.88 54.746 ;
        RECT 36.774 54.715 41.834 54.792 ;
        RECT 36.728 54.761 41.788 54.838 ;
        RECT 36.682 54.807 41.742 54.884 ;
        RECT 36.636 54.853 41.696 54.93 ;
        RECT 36.59 54.899 41.65 54.976 ;
        RECT 36.544 54.945 41.604 55.022 ;
        RECT 36.498 54.991 41.558 55.068 ;
        RECT 36.452 55.037 41.512 55.114 ;
        RECT 36.406 55.083 41.466 55.16 ;
        RECT 36.36 55.129 41.42 55.206 ;
        RECT 36.314 55.175 41.374 55.252 ;
        RECT 36.268 55.221 41.328 55.298 ;
        RECT 36.222 55.267 41.282 55.344 ;
        RECT 36.176 55.313 41.236 55.39 ;
        RECT 36.13 55.359 41.19 55.436 ;
        RECT 36.084 55.405 41.144 55.482 ;
        RECT 36.038 55.451 41.098 55.528 ;
        RECT 35.992 55.497 41.052 55.574 ;
        RECT 35.946 55.543 41.006 55.62 ;
        RECT 35.9 55.589 40.96 55.666 ;
        RECT 35.854 55.635 40.914 55.712 ;
        RECT 35.808 55.681 40.868 55.758 ;
        RECT 35.762 55.727 40.822 55.804 ;
        RECT 35.716 55.773 40.776 55.85 ;
        RECT 35.67 55.819 40.73 55.896 ;
        RECT 35.624 55.865 40.684 55.942 ;
        RECT 35.578 55.911 40.638 55.988 ;
        RECT 35.532 55.957 40.592 56.034 ;
        RECT 35.486 56.003 40.546 56.08 ;
        RECT 35.44 56.049 40.5 56.126 ;
        RECT 35.394 56.095 40.454 56.172 ;
        RECT 35.348 56.141 40.408 56.218 ;
        RECT 35.302 56.187 40.362 56.264 ;
        RECT 35.256 56.233 40.316 56.31 ;
        RECT 35.21 56.279 40.27 56.356 ;
        RECT 35.164 56.325 40.224 56.402 ;
        RECT 35.118 56.371 40.178 56.448 ;
        RECT 35.072 56.417 40.132 56.494 ;
        RECT 35.026 56.463 40.086 56.54 ;
        RECT 34.98 56.509 40.04 56.586 ;
        RECT 34.934 56.555 39.994 56.632 ;
        RECT 34.888 56.601 39.948 56.678 ;
        RECT 34.842 56.647 39.902 56.724 ;
        RECT 34.75 56.739 39.856 56.77 ;
        RECT 34.796 56.693 39.856 56.77 ;
        RECT 34.738 56.768 39.81 56.816 ;
        RECT 34.692 56.797 39.764 56.862 ;
        RECT 34.646 56.843 39.718 56.908 ;
        RECT 34.6 56.889 39.672 56.954 ;
        RECT 34.554 56.935 39.626 57 ;
        RECT 34.508 56.981 39.58 57.046 ;
        RECT 34.462 57.027 39.534 57.092 ;
        RECT 34.416 57.073 39.488 57.138 ;
        RECT 34.37 57.119 39.442 57.184 ;
        RECT 34.324 57.165 39.396 57.23 ;
        RECT 34.278 57.211 39.35 57.276 ;
        RECT 34.232 57.257 39.304 57.322 ;
        RECT 34.186 57.303 39.258 57.368 ;
        RECT 34.14 57.349 39.212 57.414 ;
        RECT 34.094 57.395 39.166 57.46 ;
        RECT 34.048 57.441 39.12 57.506 ;
        RECT 34.002 57.487 39.074 57.552 ;
        RECT 33.956 57.533 39.028 57.598 ;
        RECT 33.91 57.579 38.982 57.644 ;
        RECT 33.864 57.625 38.936 57.69 ;
        RECT 33.818 57.671 38.89 57.736 ;
        RECT 33.772 57.717 38.844 57.782 ;
        RECT 33.726 57.763 38.798 57.828 ;
        RECT 33.68 57.809 38.752 57.874 ;
        RECT 33.634 57.855 38.706 57.92 ;
        RECT 33.588 57.901 38.66 57.966 ;
        RECT 33.542 57.947 38.614 58.012 ;
        RECT 33.496 57.993 38.568 58.058 ;
        RECT 33.45 58.039 38.522 58.104 ;
        RECT 33.404 58.085 38.476 58.15 ;
        RECT 33.358 58.131 38.43 58.196 ;
        RECT 33.312 58.177 38.384 58.242 ;
        RECT 33.266 58.223 38.338 58.288 ;
        RECT 33.22 58.269 38.292 58.334 ;
        RECT 33.174 58.315 38.246 58.38 ;
        RECT 33.128 58.361 38.2 58.426 ;
        RECT 33.082 58.407 38.154 58.472 ;
        RECT 33.036 58.453 38.108 58.518 ;
        RECT 32.99 58.499 38.062 58.564 ;
        RECT 32.944 58.545 38.016 58.61 ;
        RECT 32.898 58.591 37.97 58.656 ;
        RECT 32.852 58.637 37.924 58.702 ;
        RECT 32.806 58.683 37.878 58.748 ;
        RECT 32.76 58.729 37.832 58.794 ;
        RECT 32.714 58.775 37.786 58.84 ;
        RECT 32.668 58.821 37.74 58.886 ;
        RECT 32.622 58.867 37.694 58.932 ;
        RECT 32.576 58.913 37.648 58.978 ;
        RECT 32.53 58.959 37.602 59.024 ;
        RECT 32.484 59.005 37.556 59.07 ;
        RECT 32.438 59.051 37.51 59.116 ;
        RECT 32.392 59.097 37.464 59.162 ;
        RECT 32.346 59.143 37.418 59.208 ;
        RECT 32.3 59.189 37.372 59.254 ;
        RECT 32.254 59.235 37.326 59.3 ;
        RECT 32.208 59.281 37.28 59.346 ;
        RECT 32.162 59.327 37.234 59.392 ;
        RECT 32.116 59.373 37.188 59.438 ;
        RECT 32.07 59.419 37.142 59.484 ;
        RECT 32.024 59.465 37.096 59.53 ;
        RECT 31.978 59.511 37.05 59.576 ;
        RECT 31.932 59.557 37.004 59.622 ;
        RECT 31.886 59.603 36.958 59.668 ;
        RECT 31.84 59.649 36.912 59.714 ;
        RECT 31.794 59.695 36.866 59.76 ;
        RECT 31.748 59.741 36.82 59.806 ;
        RECT 31.702 59.787 36.774 59.852 ;
        RECT 31.656 59.833 36.728 59.898 ;
        RECT 31.61 59.879 36.682 59.944 ;
        RECT 31.564 59.925 36.636 59.99 ;
        RECT 31.518 59.971 36.59 60.036 ;
        RECT 31.472 60.017 36.544 60.082 ;
        RECT 31.426 60.063 36.498 60.128 ;
        RECT 31.38 60.109 36.452 60.174 ;
        RECT 31.334 60.155 36.406 60.22 ;
        RECT 31.288 60.201 36.36 60.266 ;
        RECT 31.242 60.247 36.314 60.312 ;
        RECT 31.196 60.293 36.268 60.358 ;
        RECT 31.15 60.339 36.222 60.404 ;
        RECT 31.15 60.339 36.176 60.45 ;
        RECT 31.15 60.339 36.13 60.496 ;
        RECT 31.15 60.339 36.084 60.542 ;
        RECT 31.15 60.339 36.038 60.588 ;
        RECT 31.15 60.339 35.992 60.634 ;
        RECT 31.15 60.339 35.946 60.68 ;
        RECT 31.15 60.339 35.9 60.726 ;
        RECT 31.15 60.339 35.854 60.772 ;
        RECT 31.15 60.339 35.808 60.818 ;
        RECT 31.15 60.339 35.762 60.864 ;
        RECT 31.15 60.339 35.716 60.91 ;
        RECT 31.15 60.339 35.67 60.956 ;
        RECT 31.15 60.339 35.624 61.002 ;
        RECT 31.15 60.339 35.578 61.048 ;
        RECT 31.15 60.339 35.532 61.094 ;
        RECT 31.15 60.339 35.486 61.14 ;
        RECT 31.15 60.339 35.44 61.186 ;
        RECT 31.15 60.339 35.394 61.232 ;
        RECT 31.15 60.339 35.348 61.278 ;
        RECT 31.15 60.339 35.302 61.324 ;
        RECT 31.15 60.339 35.256 61.37 ;
        RECT 31.15 60.339 35.21 61.416 ;
        RECT 31.15 60.339 35.164 61.462 ;
        RECT 31.15 60.339 35.118 61.508 ;
        RECT 31.15 60.339 35.072 61.554 ;
        RECT 31.15 60.339 35.026 61.6 ;
        RECT 31.15 60.339 34.98 61.646 ;
        RECT 31.15 60.339 34.934 61.692 ;
        RECT 31.15 60.339 34.888 61.738 ;
        RECT 31.15 60.339 34.842 61.784 ;
        RECT 31.15 60.339 34.796 61.83 ;
        RECT 31.15 60.339 34.75 80 ;
    END
    PORT
      LAYER IB ;
        RECT 18.526 53.019 23.586 53.096 ;
        RECT 18.48 53.065 23.54 53.142 ;
        RECT 18.434 53.111 23.494 53.188 ;
        RECT 18.388 53.157 23.448 53.234 ;
        RECT 18.342 53.203 23.402 53.28 ;
        RECT 18.296 53.249 23.356 53.326 ;
        RECT 18.25 53.295 23.31 53.372 ;
        RECT 18.204 53.341 23.264 53.418 ;
        RECT 18.158 53.387 23.218 53.464 ;
        RECT 18.112 53.433 23.172 53.51 ;
        RECT 18.066 53.479 23.126 53.556 ;
        RECT 18.02 53.525 23.08 53.602 ;
        RECT 17.974 53.571 23.034 53.648 ;
        RECT 17.928 53.617 22.988 53.694 ;
        RECT 17.882 53.663 22.942 53.74 ;
        RECT 17.836 53.709 22.896 53.786 ;
        RECT 17.79 53.755 22.85 53.832 ;
        RECT 17.744 53.801 22.804 53.878 ;
        RECT 17.698 53.847 22.758 53.924 ;
        RECT 17.652 53.893 22.712 53.97 ;
        RECT 17.606 53.939 22.666 54.016 ;
        RECT 17.56 53.985 22.62 54.062 ;
        RECT 17.514 54.031 22.574 54.108 ;
        RECT 17.468 54.077 22.528 54.154 ;
        RECT 17.422 54.123 22.482 54.2 ;
        RECT 17.376 54.169 22.436 54.246 ;
        RECT 17.33 54.215 22.39 54.292 ;
        RECT 17.284 54.261 22.344 54.338 ;
        RECT 17.238 54.307 22.298 54.384 ;
        RECT 17.192 54.353 22.252 54.43 ;
        RECT 17.146 54.399 22.206 54.476 ;
        RECT 17.1 54.445 22.16 54.522 ;
        RECT 17.054 54.491 22.114 54.568 ;
        RECT 17.008 54.537 22.068 54.614 ;
        RECT 16.962 54.583 22.022 54.66 ;
        RECT 16.916 54.629 21.976 54.706 ;
        RECT 16.87 54.675 21.93 54.752 ;
        RECT 16.824 54.721 21.884 54.798 ;
        RECT 16.778 54.767 21.838 54.844 ;
        RECT 16.732 54.813 21.792 54.89 ;
        RECT 16.686 54.859 21.746 54.936 ;
        RECT 16.64 54.905 21.7 54.982 ;
        RECT 16.594 54.951 21.654 55.028 ;
        RECT 16.548 54.997 21.608 55.074 ;
        RECT 16.502 55.043 21.562 55.12 ;
        RECT 16.456 55.089 21.516 55.166 ;
        RECT 16.41 55.135 21.47 55.212 ;
        RECT 16.364 55.181 21.424 55.258 ;
        RECT 16.318 55.227 21.378 55.304 ;
        RECT 16.272 55.273 21.332 55.35 ;
        RECT 16.226 55.319 21.286 55.396 ;
        RECT 16.18 55.365 21.24 55.442 ;
        RECT 16.134 55.411 21.194 55.488 ;
        RECT 16.088 55.457 21.148 55.534 ;
        RECT 16.042 55.503 21.102 55.58 ;
        RECT 15.95 55.595 21.056 55.626 ;
        RECT 15.996 55.549 21.056 55.626 ;
        RECT 15.938 55.624 21.01 55.672 ;
        RECT 15.892 55.653 20.964 55.718 ;
        RECT 15.846 55.699 20.918 55.764 ;
        RECT 15.8 55.745 20.872 55.81 ;
        RECT 15.754 55.791 20.826 55.856 ;
        RECT 15.708 55.837 20.78 55.902 ;
        RECT 15.662 55.883 20.734 55.948 ;
        RECT 15.616 55.929 20.688 55.994 ;
        RECT 15.57 55.975 20.642 56.04 ;
        RECT 15.524 56.021 20.596 56.086 ;
        RECT 15.478 56.067 20.55 56.132 ;
        RECT 15.432 56.113 20.504 56.178 ;
        RECT 15.386 56.159 20.458 56.224 ;
        RECT 15.34 56.205 20.412 56.27 ;
        RECT 15.294 56.251 20.366 56.316 ;
        RECT 15.248 56.297 20.32 56.362 ;
        RECT 15.202 56.343 20.274 56.408 ;
        RECT 15.156 56.389 20.228 56.454 ;
        RECT 15.11 56.435 20.182 56.5 ;
        RECT 15.064 56.481 20.136 56.546 ;
        RECT 15.018 56.527 20.09 56.592 ;
        RECT 14.972 56.573 20.044 56.638 ;
        RECT 14.926 56.619 19.998 56.684 ;
        RECT 14.88 56.665 19.952 56.73 ;
        RECT 14.834 56.711 19.906 56.776 ;
        RECT 14.788 56.757 19.86 56.822 ;
        RECT 14.742 56.803 19.814 56.868 ;
        RECT 14.696 56.849 19.768 56.914 ;
        RECT 14.65 56.895 19.722 56.96 ;
        RECT 14.604 56.941 19.676 57.006 ;
        RECT 14.558 56.987 19.63 57.052 ;
        RECT 14.512 57.033 19.584 57.098 ;
        RECT 14.466 57.079 19.538 57.144 ;
        RECT 14.42 57.125 19.492 57.19 ;
        RECT 14.374 57.171 19.446 57.236 ;
        RECT 14.328 57.217 19.4 57.282 ;
        RECT 14.282 57.263 19.354 57.328 ;
        RECT 14.236 57.309 19.308 57.374 ;
        RECT 14.19 57.355 19.262 57.42 ;
        RECT 14.144 57.401 19.216 57.466 ;
        RECT 14.098 57.447 19.17 57.512 ;
        RECT 14.052 57.493 19.124 57.558 ;
        RECT 14.006 57.539 19.078 57.604 ;
        RECT 13.96 57.585 19.032 57.65 ;
        RECT 13.914 57.631 18.986 57.696 ;
        RECT 13.868 57.677 18.94 57.742 ;
        RECT 13.822 57.723 18.894 57.788 ;
        RECT 13.776 57.769 18.848 57.834 ;
        RECT 13.73 57.815 18.802 57.88 ;
        RECT 13.684 57.861 18.756 57.926 ;
        RECT 13.638 57.907 18.71 57.972 ;
        RECT 13.592 57.953 18.664 58.018 ;
        RECT 13.546 57.999 18.618 58.064 ;
        RECT 13.5 58.045 18.572 58.11 ;
        RECT 13.454 58.091 18.526 58.156 ;
        RECT 13.408 58.137 18.48 58.202 ;
        RECT 13.362 58.183 18.434 58.248 ;
        RECT 13.316 58.229 18.388 58.294 ;
        RECT 13.27 58.275 18.342 58.34 ;
        RECT 13.224 58.321 18.296 58.386 ;
        RECT 13.178 58.367 18.25 58.432 ;
        RECT 13.132 58.413 18.204 58.478 ;
        RECT 13.086 58.459 18.158 58.524 ;
        RECT 13.04 58.505 18.112 58.57 ;
        RECT 12.994 58.551 18.066 58.616 ;
        RECT 12.948 58.597 18.02 58.662 ;
        RECT 12.902 58.643 17.974 58.708 ;
        RECT 12.856 58.689 17.928 58.754 ;
        RECT 12.81 58.735 17.882 58.8 ;
        RECT 12.764 58.781 17.836 58.846 ;
        RECT 12.718 58.827 17.79 58.892 ;
        RECT 12.672 58.873 17.744 58.938 ;
        RECT 12.626 58.919 17.698 58.984 ;
        RECT 12.58 58.965 17.652 59.03 ;
        RECT 12.534 59.011 17.606 59.076 ;
        RECT 12.488 59.057 17.56 59.122 ;
        RECT 12.442 59.103 17.514 59.168 ;
        RECT 12.396 59.149 17.468 59.214 ;
        RECT 12.35 59.195 17.422 59.26 ;
        RECT 12.35 59.195 17.376 59.306 ;
        RECT 12.35 59.195 17.33 59.352 ;
        RECT 12.35 59.195 17.284 59.398 ;
        RECT 12.35 59.195 17.238 59.444 ;
        RECT 12.35 59.195 17.192 59.49 ;
        RECT 12.35 59.195 17.146 59.536 ;
        RECT 12.35 59.195 17.1 59.582 ;
        RECT 12.35 59.195 17.054 59.628 ;
        RECT 12.35 59.195 17.008 59.674 ;
        RECT 12.35 59.195 16.962 59.72 ;
        RECT 12.35 59.195 16.916 59.766 ;
        RECT 12.35 59.195 16.87 59.812 ;
        RECT 12.35 59.195 16.824 59.858 ;
        RECT 12.35 59.195 16.778 59.904 ;
        RECT 12.35 59.195 16.732 59.95 ;
        RECT 12.35 59.195 16.686 59.996 ;
        RECT 12.35 59.195 16.64 60.042 ;
        RECT 12.35 59.195 16.594 60.088 ;
        RECT 12.35 59.195 16.548 60.134 ;
        RECT 12.35 59.195 16.502 60.18 ;
        RECT 12.35 59.195 16.456 60.226 ;
        RECT 12.35 59.195 16.41 60.272 ;
        RECT 12.35 59.195 16.364 60.318 ;
        RECT 12.35 59.195 16.318 60.364 ;
        RECT 12.35 59.195 16.272 60.41 ;
        RECT 12.35 59.195 16.226 60.456 ;
        RECT 12.35 59.195 16.18 60.502 ;
        RECT 12.35 59.195 16.134 60.548 ;
        RECT 12.35 59.195 16.088 60.594 ;
        RECT 12.35 59.195 16.042 60.64 ;
        RECT 12.35 59.195 15.996 60.686 ;
        RECT 12.35 59.195 15.95 80 ;
        RECT 59.218 12.35 80 15.95 ;
        RECT 55.602 15.943 60.709 15.96 ;
        RECT 54.176 17.369 59.264 17.418 ;
        RECT 59.19 12.364 59.218 17.455 ;
        RECT 54.13 17.415 59.19 17.492 ;
        RECT 54.222 17.323 59.31 17.372 ;
        RECT 59.144 12.401 59.19 17.492 ;
        RECT 54.084 17.461 59.144 17.538 ;
        RECT 54.268 17.277 59.356 17.326 ;
        RECT 59.098 12.447 59.144 17.538 ;
        RECT 54.038 17.507 59.098 17.584 ;
        RECT 54.314 17.231 59.402 17.28 ;
        RECT 59.052 12.493 59.098 17.584 ;
        RECT 53.992 17.553 59.052 17.63 ;
        RECT 54.36 17.185 59.448 17.234 ;
        RECT 59.006 12.539 59.052 17.63 ;
        RECT 53.946 17.599 59.006 17.676 ;
        RECT 54.406 17.139 59.494 17.188 ;
        RECT 58.96 12.585 59.006 17.676 ;
        RECT 53.9 17.645 58.96 17.722 ;
        RECT 54.452 17.093 59.54 17.142 ;
        RECT 58.914 12.631 58.96 17.722 ;
        RECT 53.854 17.691 58.914 17.768 ;
        RECT 54.498 17.047 59.586 17.096 ;
        RECT 58.868 12.677 58.914 17.768 ;
        RECT 53.808 17.737 58.868 17.814 ;
        RECT 54.544 17.001 59.632 17.05 ;
        RECT 58.822 12.723 58.868 17.814 ;
        RECT 53.762 17.783 58.822 17.86 ;
        RECT 54.59 16.955 59.678 17.004 ;
        RECT 58.776 12.769 58.822 17.86 ;
        RECT 53.716 17.829 58.776 17.906 ;
        RECT 54.636 16.909 59.724 16.958 ;
        RECT 58.73 12.815 58.776 17.906 ;
        RECT 53.67 17.875 58.73 17.952 ;
        RECT 54.682 16.863 59.77 16.912 ;
        RECT 58.684 12.861 58.73 17.952 ;
        RECT 53.624 17.921 58.684 17.998 ;
        RECT 54.728 16.817 59.816 16.866 ;
        RECT 58.638 12.907 58.684 17.998 ;
        RECT 53.578 17.967 58.638 18.044 ;
        RECT 54.774 16.771 59.862 16.82 ;
        RECT 58.592 12.953 58.638 18.044 ;
        RECT 53.532 18.013 58.592 18.09 ;
        RECT 54.82 16.725 59.908 16.774 ;
        RECT 58.546 12.999 58.592 18.09 ;
        RECT 53.486 18.059 58.546 18.136 ;
        RECT 54.866 16.679 59.954 16.728 ;
        RECT 58.5 13.045 58.546 18.136 ;
        RECT 53.44 18.105 58.5 18.182 ;
        RECT 54.912 16.633 60 16.682 ;
        RECT 58.454 13.091 58.5 18.182 ;
        RECT 53.394 18.151 58.454 18.228 ;
        RECT 54.958 16.587 60.046 16.636 ;
        RECT 58.408 13.137 58.454 18.228 ;
        RECT 53.348 18.197 58.408 18.274 ;
        RECT 55.004 16.541 60.092 16.59 ;
        RECT 58.362 13.183 58.408 18.274 ;
        RECT 53.302 18.243 58.362 18.32 ;
        RECT 55.05 16.495 60.138 16.544 ;
        RECT 58.316 13.229 58.362 18.32 ;
        RECT 53.256 18.289 58.316 18.366 ;
        RECT 55.096 16.449 60.184 16.498 ;
        RECT 58.27 13.275 58.316 18.366 ;
        RECT 53.21 18.335 58.27 18.412 ;
        RECT 55.142 16.403 60.23 16.452 ;
        RECT 58.224 13.321 58.27 18.412 ;
        RECT 53.164 18.381 58.224 18.458 ;
        RECT 55.188 16.357 60.276 16.406 ;
        RECT 58.178 13.367 58.224 18.458 ;
        RECT 53.118 18.427 58.178 18.504 ;
        RECT 55.234 16.311 60.322 16.36 ;
        RECT 58.132 13.413 58.178 18.504 ;
        RECT 53.072 18.473 58.132 18.55 ;
        RECT 55.28 16.265 60.368 16.314 ;
        RECT 58.086 13.459 58.132 18.55 ;
        RECT 53.026 18.519 58.086 18.596 ;
        RECT 55.326 16.219 60.414 16.268 ;
        RECT 58.04 13.505 58.086 18.596 ;
        RECT 52.98 18.565 58.04 18.642 ;
        RECT 55.372 16.173 60.46 16.222 ;
        RECT 57.994 13.551 58.04 18.642 ;
        RECT 52.934 18.611 57.994 18.688 ;
        RECT 55.418 16.127 60.506 16.176 ;
        RECT 57.948 13.597 57.994 18.688 ;
        RECT 52.888 18.657 57.948 18.734 ;
        RECT 55.464 16.081 60.552 16.13 ;
        RECT 57.902 13.643 57.948 18.734 ;
        RECT 52.842 18.703 57.902 18.78 ;
        RECT 55.51 16.035 60.598 16.084 ;
        RECT 57.856 13.689 57.902 18.78 ;
        RECT 52.796 18.749 57.856 18.826 ;
        RECT 55.556 15.989 60.644 16.038 ;
        RECT 57.81 13.735 57.856 18.826 ;
        RECT 52.75 18.795 57.81 18.872 ;
        RECT 55.602 15.943 60.69 15.992 ;
        RECT 57.764 13.781 57.81 18.872 ;
        RECT 52.704 18.841 57.764 18.918 ;
        RECT 55.648 15.897 80 15.95 ;
        RECT 57.718 13.827 57.764 18.918 ;
        RECT 52.658 18.887 57.718 18.964 ;
        RECT 55.694 15.851 80 15.95 ;
        RECT 57.672 13.873 57.718 18.964 ;
        RECT 52.612 18.933 57.672 19.01 ;
        RECT 55.74 15.805 80 15.95 ;
        RECT 57.626 13.919 57.672 19.01 ;
        RECT 52.566 18.979 57.626 19.056 ;
        RECT 55.786 15.759 80 15.95 ;
        RECT 57.58 13.965 57.626 19.056 ;
        RECT 52.52 19.025 57.58 19.102 ;
        RECT 55.832 15.713 80 15.95 ;
        RECT 57.534 14.011 57.58 19.102 ;
        RECT 52.474 19.071 57.534 19.148 ;
        RECT 55.878 15.667 80 15.95 ;
        RECT 57.488 14.057 57.534 19.148 ;
        RECT 52.428 19.117 57.488 19.194 ;
        RECT 55.924 15.621 80 15.95 ;
        RECT 57.442 14.103 57.488 19.194 ;
        RECT 52.382 19.163 57.442 19.24 ;
        RECT 55.97 15.575 80 15.95 ;
        RECT 57.396 14.149 57.442 19.24 ;
        RECT 52.336 19.209 57.396 19.286 ;
        RECT 56.016 15.529 80 15.95 ;
        RECT 57.35 14.195 57.396 19.286 ;
        RECT 52.29 19.255 57.35 19.332 ;
        RECT 56.062 15.483 80 15.95 ;
        RECT 57.304 14.241 57.35 19.332 ;
        RECT 52.244 19.301 57.304 19.378 ;
        RECT 56.108 15.437 80 15.95 ;
        RECT 57.258 14.287 57.304 19.378 ;
        RECT 52.198 19.347 57.258 19.424 ;
        RECT 56.154 15.391 80 15.95 ;
        RECT 57.212 14.333 57.258 19.424 ;
        RECT 52.152 19.393 57.212 19.47 ;
        RECT 56.2 15.345 80 15.95 ;
        RECT 57.166 14.379 57.212 19.47 ;
        RECT 52.106 19.439 57.166 19.516 ;
        RECT 56.246 15.299 80 15.95 ;
        RECT 57.12 14.425 57.166 19.516 ;
        RECT 52.06 19.485 57.12 19.562 ;
        RECT 56.292 15.253 80 15.95 ;
        RECT 57.074 14.471 57.12 19.562 ;
        RECT 52.014 19.531 57.074 19.608 ;
        RECT 56.338 15.207 80 15.95 ;
        RECT 57.028 14.517 57.074 19.608 ;
        RECT 51.968 19.577 57.028 19.654 ;
        RECT 56.384 15.161 80 15.95 ;
        RECT 56.982 14.563 57.028 19.654 ;
        RECT 51.922 19.623 56.982 19.7 ;
        RECT 56.43 15.115 80 15.95 ;
        RECT 56.936 14.609 56.982 19.7 ;
        RECT 51.876 19.669 56.936 19.746 ;
        RECT 56.476 15.069 80 15.95 ;
        RECT 56.89 14.655 56.936 19.746 ;
        RECT 51.83 19.715 56.89 19.792 ;
        RECT 56.522 15.023 80 15.95 ;
        RECT 56.844 14.701 56.89 19.792 ;
        RECT 51.784 19.761 56.844 19.838 ;
        RECT 56.568 14.977 80 15.95 ;
        RECT 56.798 14.747 56.844 19.838 ;
        RECT 51.738 19.807 56.798 19.884 ;
        RECT 56.614 14.931 80 15.95 ;
        RECT 56.752 14.793 56.798 19.884 ;
        RECT 51.692 19.853 56.752 19.93 ;
        RECT 56.66 14.885 80 15.95 ;
        RECT 56.706 14.839 56.752 19.93 ;
        RECT 51.646 19.899 56.706 19.976 ;
        RECT 51.6 19.945 56.66 20.022 ;
        RECT 51.554 19.991 56.614 20.068 ;
        RECT 51.508 20.037 56.568 20.114 ;
        RECT 51.462 20.083 56.522 20.16 ;
        RECT 51.416 20.129 56.476 20.206 ;
        RECT 51.37 20.175 56.43 20.252 ;
        RECT 51.324 20.221 56.384 20.298 ;
        RECT 51.278 20.267 56.338 20.344 ;
        RECT 51.232 20.313 56.292 20.39 ;
        RECT 51.186 20.359 56.246 20.436 ;
        RECT 51.14 20.405 56.2 20.482 ;
        RECT 51.094 20.451 56.154 20.528 ;
        RECT 51.048 20.497 56.108 20.574 ;
        RECT 51.002 20.543 56.062 20.62 ;
        RECT 50.956 20.589 56.016 20.666 ;
        RECT 50.91 20.635 55.97 20.712 ;
        RECT 50.864 20.681 55.924 20.758 ;
        RECT 50.818 20.727 55.878 20.804 ;
        RECT 50.772 20.773 55.832 20.85 ;
        RECT 50.726 20.819 55.786 20.896 ;
        RECT 50.68 20.865 55.74 20.942 ;
        RECT 50.634 20.911 55.694 20.988 ;
        RECT 50.588 20.957 55.648 21.034 ;
        RECT 50.542 21.003 55.602 21.08 ;
        RECT 50.496 21.049 55.556 21.126 ;
        RECT 50.45 21.095 55.51 21.172 ;
        RECT 50.404 21.141 55.464 21.218 ;
        RECT 50.358 21.187 55.418 21.264 ;
        RECT 50.312 21.233 55.372 21.31 ;
        RECT 50.266 21.279 55.326 21.356 ;
        RECT 50.22 21.325 55.28 21.402 ;
        RECT 50.174 21.371 55.234 21.448 ;
        RECT 50.128 21.417 55.188 21.494 ;
        RECT 50.082 21.463 55.142 21.54 ;
        RECT 50.036 21.509 55.096 21.586 ;
        RECT 49.99 21.555 55.05 21.632 ;
        RECT 49.944 21.601 55.004 21.678 ;
        RECT 49.898 21.647 54.958 21.724 ;
        RECT 49.852 21.693 54.912 21.77 ;
        RECT 49.806 21.739 54.866 21.816 ;
        RECT 49.76 21.785 54.82 21.862 ;
        RECT 49.714 21.831 54.774 21.908 ;
        RECT 49.668 21.877 54.728 21.954 ;
        RECT 49.622 21.923 54.682 22 ;
        RECT 49.576 21.969 54.636 22.046 ;
        RECT 49.53 22.015 54.59 22.092 ;
        RECT 49.484 22.061 54.544 22.138 ;
        RECT 49.438 22.107 54.498 22.184 ;
        RECT 49.392 22.153 54.452 22.23 ;
        RECT 49.346 22.199 54.406 22.276 ;
        RECT 49.3 22.245 54.36 22.322 ;
        RECT 49.254 22.291 54.314 22.368 ;
        RECT 49.208 22.337 54.268 22.414 ;
        RECT 49.162 22.383 54.222 22.46 ;
        RECT 49.116 22.429 54.176 22.506 ;
        RECT 49.07 22.475 54.13 22.552 ;
        RECT 49.024 22.521 54.084 22.598 ;
        RECT 48.978 22.567 54.038 22.644 ;
        RECT 48.932 22.613 53.992 22.69 ;
        RECT 48.886 22.659 53.946 22.736 ;
        RECT 48.84 22.705 53.9 22.782 ;
        RECT 48.794 22.751 53.854 22.828 ;
        RECT 48.748 22.797 53.808 22.874 ;
        RECT 48.702 22.843 53.762 22.92 ;
        RECT 48.656 22.889 53.716 22.966 ;
        RECT 48.61 22.935 53.67 23.012 ;
        RECT 48.564 22.981 53.624 23.058 ;
        RECT 48.518 23.027 53.578 23.104 ;
        RECT 48.472 23.073 53.532 23.15 ;
        RECT 48.426 23.119 53.486 23.196 ;
        RECT 48.38 23.165 53.44 23.242 ;
        RECT 48.334 23.211 53.394 23.288 ;
        RECT 48.288 23.257 53.348 23.334 ;
        RECT 48.242 23.303 53.302 23.38 ;
        RECT 48.196 23.349 53.256 23.426 ;
        RECT 48.15 23.395 53.21 23.472 ;
        RECT 48.104 23.441 53.164 23.518 ;
        RECT 48.058 23.487 53.118 23.564 ;
        RECT 48.012 23.533 53.072 23.61 ;
        RECT 47.966 23.579 53.026 23.656 ;
        RECT 47.92 23.625 52.98 23.702 ;
        RECT 47.874 23.671 52.934 23.748 ;
        RECT 47.828 23.717 52.888 23.794 ;
        RECT 47.782 23.763 52.842 23.84 ;
        RECT 47.736 23.809 52.796 23.886 ;
        RECT 47.69 23.855 52.75 23.932 ;
        RECT 47.644 23.901 52.704 23.978 ;
        RECT 47.598 23.947 52.658 24.024 ;
        RECT 47.552 23.993 52.612 24.07 ;
        RECT 47.506 24.039 52.566 24.116 ;
        RECT 47.46 24.085 52.52 24.162 ;
        RECT 47.414 24.131 52.474 24.208 ;
        RECT 47.368 24.177 52.428 24.254 ;
        RECT 47.322 24.223 52.382 24.3 ;
        RECT 47.276 24.269 52.336 24.346 ;
        RECT 47.23 24.315 52.29 24.392 ;
        RECT 47.184 24.361 52.244 24.438 ;
        RECT 47.138 24.407 52.198 24.484 ;
        RECT 47.092 24.453 52.152 24.53 ;
        RECT 47.046 24.499 52.106 24.576 ;
        RECT 47 24.545 52.06 24.622 ;
        RECT 46.954 24.591 52.014 24.668 ;
        RECT 46.908 24.637 51.968 24.714 ;
        RECT 46.862 24.683 51.922 24.76 ;
        RECT 46.816 24.729 51.876 24.806 ;
        RECT 46.77 24.775 51.83 24.852 ;
        RECT 46.724 24.821 51.784 24.898 ;
        RECT 46.678 24.867 51.738 24.944 ;
        RECT 46.632 24.913 51.692 24.99 ;
        RECT 46.586 24.959 51.646 25.036 ;
        RECT 46.54 25.005 51.6 25.082 ;
        RECT 46.494 25.051 51.554 25.128 ;
        RECT 46.448 25.097 51.508 25.174 ;
        RECT 46.402 25.143 51.462 25.22 ;
        RECT 46.356 25.189 51.416 25.266 ;
        RECT 46.31 25.235 51.37 25.312 ;
        RECT 46.264 25.281 51.324 25.358 ;
        RECT 46.218 25.327 51.278 25.404 ;
        RECT 46.172 25.373 51.232 25.45 ;
        RECT 46.126 25.419 51.186 25.496 ;
        RECT 46.08 25.465 51.14 25.542 ;
        RECT 46.034 25.511 51.094 25.588 ;
        RECT 45.988 25.557 51.048 25.634 ;
        RECT 45.942 25.603 51.002 25.68 ;
        RECT 45.896 25.649 50.956 25.726 ;
        RECT 45.85 25.695 50.91 25.772 ;
        RECT 45.804 25.741 50.864 25.818 ;
        RECT 45.758 25.787 50.818 25.864 ;
        RECT 45.712 25.833 50.772 25.91 ;
        RECT 45.666 25.879 50.726 25.956 ;
        RECT 45.62 25.925 50.68 26.002 ;
        RECT 45.574 25.971 50.634 26.048 ;
        RECT 45.528 26.017 50.588 26.094 ;
        RECT 45.482 26.063 50.542 26.14 ;
        RECT 45.436 26.109 50.496 26.186 ;
        RECT 45.39 26.155 50.45 26.232 ;
        RECT 45.344 26.201 50.404 26.278 ;
        RECT 45.298 26.247 50.358 26.324 ;
        RECT 45.252 26.293 50.312 26.37 ;
        RECT 45.206 26.339 50.266 26.416 ;
        RECT 45.16 26.385 50.22 26.462 ;
        RECT 45.114 26.431 50.174 26.508 ;
        RECT 45.068 26.477 50.128 26.554 ;
        RECT 45.022 26.523 50.082 26.6 ;
        RECT 44.976 26.569 50.036 26.646 ;
        RECT 44.93 26.615 49.99 26.692 ;
        RECT 44.884 26.661 49.944 26.738 ;
        RECT 44.838 26.707 49.898 26.784 ;
        RECT 44.792 26.753 49.852 26.83 ;
        RECT 44.746 26.799 49.806 26.876 ;
        RECT 44.7 26.845 49.76 26.922 ;
        RECT 44.654 26.891 49.714 26.968 ;
        RECT 44.608 26.937 49.668 27.014 ;
        RECT 44.562 26.983 49.622 27.06 ;
        RECT 44.516 27.029 49.576 27.106 ;
        RECT 44.47 27.075 49.53 27.152 ;
        RECT 44.424 27.121 49.484 27.198 ;
        RECT 44.378 27.167 49.438 27.244 ;
        RECT 44.332 27.213 49.392 27.29 ;
        RECT 44.286 27.259 49.346 27.336 ;
        RECT 44.24 27.305 49.3 27.382 ;
        RECT 44.194 27.351 49.254 27.428 ;
        RECT 44.148 27.397 49.208 27.474 ;
        RECT 44.102 27.443 49.162 27.52 ;
        RECT 44.056 27.489 49.116 27.566 ;
        RECT 44.01 27.535 49.07 27.612 ;
        RECT 43.964 27.581 49.024 27.658 ;
        RECT 43.918 27.627 48.978 27.704 ;
        RECT 43.872 27.673 48.932 27.75 ;
        RECT 43.826 27.719 48.886 27.796 ;
        RECT 43.78 27.765 48.84 27.842 ;
        RECT 43.734 27.811 48.794 27.888 ;
        RECT 43.688 27.857 48.748 27.934 ;
        RECT 43.642 27.903 48.702 27.98 ;
        RECT 43.596 27.949 48.656 28.026 ;
        RECT 43.55 27.995 48.61 28.072 ;
        RECT 43.504 28.041 48.564 28.118 ;
        RECT 43.458 28.087 48.518 28.164 ;
        RECT 43.412 28.133 48.472 28.21 ;
        RECT 43.366 28.179 48.426 28.256 ;
        RECT 43.32 28.225 48.38 28.302 ;
        RECT 43.274 28.271 48.334 28.348 ;
        RECT 43.228 28.317 48.288 28.394 ;
        RECT 43.182 28.363 48.242 28.44 ;
        RECT 43.136 28.409 48.196 28.486 ;
        RECT 43.09 28.455 48.15 28.532 ;
        RECT 43.044 28.501 48.104 28.578 ;
        RECT 42.998 28.547 48.058 28.624 ;
        RECT 42.952 28.593 48.012 28.67 ;
        RECT 42.906 28.639 47.966 28.716 ;
        RECT 42.86 28.685 47.92 28.762 ;
        RECT 42.814 28.731 47.874 28.808 ;
        RECT 42.768 28.777 47.828 28.854 ;
        RECT 42.722 28.823 47.782 28.9 ;
        RECT 42.676 28.869 47.736 28.946 ;
        RECT 42.63 28.915 47.69 28.992 ;
        RECT 42.584 28.961 47.644 29.038 ;
        RECT 42.538 29.007 47.598 29.084 ;
        RECT 42.492 29.053 47.552 29.13 ;
        RECT 42.446 29.099 47.506 29.176 ;
        RECT 42.4 29.145 47.46 29.222 ;
        RECT 42.354 29.191 47.414 29.268 ;
        RECT 42.308 29.237 47.368 29.314 ;
        RECT 42.262 29.283 47.322 29.36 ;
        RECT 42.216 29.329 47.276 29.406 ;
        RECT 42.17 29.375 47.23 29.452 ;
        RECT 42.124 29.421 47.184 29.498 ;
        RECT 42.078 29.467 47.138 29.544 ;
        RECT 42.032 29.513 47.092 29.59 ;
        RECT 41.986 29.559 47.046 29.636 ;
        RECT 41.94 29.605 47 29.682 ;
        RECT 41.894 29.651 46.954 29.728 ;
        RECT 41.848 29.697 46.908 29.774 ;
        RECT 41.802 29.743 46.862 29.82 ;
        RECT 41.756 29.789 46.816 29.866 ;
        RECT 41.71 29.835 46.77 29.912 ;
        RECT 41.664 29.881 46.724 29.958 ;
        RECT 41.618 29.927 46.678 30.004 ;
        RECT 41.572 29.973 46.632 30.05 ;
        RECT 41.526 30.019 46.586 30.096 ;
        RECT 41.48 30.065 46.54 30.142 ;
        RECT 41.434 30.111 46.494 30.188 ;
        RECT 41.388 30.157 46.448 30.234 ;
        RECT 41.342 30.203 46.402 30.28 ;
        RECT 41.296 30.249 46.356 30.326 ;
        RECT 41.25 30.295 46.31 30.372 ;
        RECT 41.204 30.341 46.264 30.418 ;
        RECT 41.158 30.387 46.218 30.464 ;
        RECT 41.112 30.433 46.172 30.51 ;
        RECT 41.066 30.479 46.126 30.556 ;
        RECT 41.02 30.525 46.08 30.602 ;
        RECT 40.974 30.571 46.034 30.648 ;
        RECT 40.928 30.617 45.988 30.694 ;
        RECT 40.882 30.663 45.942 30.74 ;
        RECT 40.836 30.709 45.896 30.786 ;
        RECT 40.79 30.755 45.85 30.832 ;
        RECT 40.744 30.801 45.804 30.878 ;
        RECT 40.698 30.847 45.758 30.924 ;
        RECT 40.652 30.893 45.712 30.97 ;
        RECT 40.606 30.939 45.666 31.016 ;
        RECT 40.56 30.985 45.62 31.062 ;
        RECT 40.514 31.031 45.574 31.108 ;
        RECT 40.468 31.077 45.528 31.154 ;
        RECT 40.422 31.123 45.482 31.2 ;
        RECT 40.376 31.169 45.436 31.246 ;
        RECT 40.33 31.215 45.39 31.292 ;
        RECT 40.284 31.261 45.344 31.338 ;
        RECT 40.238 31.307 45.298 31.384 ;
        RECT 40.192 31.353 45.252 31.43 ;
        RECT 40.146 31.399 45.206 31.476 ;
        RECT 40.1 31.445 45.16 31.522 ;
        RECT 40.054 31.491 45.114 31.568 ;
        RECT 40.008 31.537 45.068 31.614 ;
        RECT 39.962 31.583 45.022 31.66 ;
        RECT 39.916 31.629 44.976 31.706 ;
        RECT 39.87 31.675 44.93 31.752 ;
        RECT 39.824 31.721 44.884 31.798 ;
        RECT 39.778 31.767 44.838 31.844 ;
        RECT 39.732 31.813 44.792 31.89 ;
        RECT 39.686 31.859 44.746 31.936 ;
        RECT 39.64 31.905 44.7 31.982 ;
        RECT 39.594 31.951 44.654 32.028 ;
        RECT 39.548 31.997 44.608 32.074 ;
        RECT 39.502 32.043 44.562 32.12 ;
        RECT 39.456 32.089 44.516 32.166 ;
        RECT 39.41 32.135 44.47 32.212 ;
        RECT 39.364 32.181 44.424 32.258 ;
        RECT 39.318 32.227 44.378 32.304 ;
        RECT 39.272 32.273 44.332 32.35 ;
        RECT 39.226 32.319 44.286 32.396 ;
        RECT 39.18 32.365 44.24 32.442 ;
        RECT 39.134 32.411 44.194 32.488 ;
        RECT 39.088 32.457 44.148 32.534 ;
        RECT 39.042 32.503 44.102 32.58 ;
        RECT 38.996 32.549 44.056 32.626 ;
        RECT 38.95 32.595 44.01 32.672 ;
        RECT 38.904 32.641 43.964 32.718 ;
        RECT 38.858 32.687 43.918 32.764 ;
        RECT 38.812 32.733 43.872 32.81 ;
        RECT 38.766 32.779 43.826 32.856 ;
        RECT 38.72 32.825 43.78 32.902 ;
        RECT 38.674 32.871 43.734 32.948 ;
        RECT 38.628 32.917 43.688 32.994 ;
        RECT 38.582 32.963 43.642 33.04 ;
        RECT 38.536 33.009 43.596 33.086 ;
        RECT 38.49 33.055 43.55 33.132 ;
        RECT 38.444 33.101 43.504 33.178 ;
        RECT 38.398 33.147 43.458 33.224 ;
        RECT 38.352 33.193 43.412 33.27 ;
        RECT 38.306 33.239 43.366 33.316 ;
        RECT 38.26 33.285 43.32 33.362 ;
        RECT 38.214 33.331 43.274 33.408 ;
        RECT 38.168 33.377 43.228 33.454 ;
        RECT 38.122 33.423 43.182 33.5 ;
        RECT 38.076 33.469 43.136 33.546 ;
        RECT 38.03 33.515 43.09 33.592 ;
        RECT 37.984 33.561 43.044 33.638 ;
        RECT 37.938 33.607 42.998 33.684 ;
        RECT 37.892 33.653 42.952 33.73 ;
        RECT 37.846 33.699 42.906 33.776 ;
        RECT 37.8 33.745 42.86 33.822 ;
        RECT 37.754 33.791 42.814 33.868 ;
        RECT 37.708 33.837 42.768 33.914 ;
        RECT 37.662 33.883 42.722 33.96 ;
        RECT 37.616 33.929 42.676 34.006 ;
        RECT 37.57 33.975 42.63 34.052 ;
        RECT 37.524 34.021 42.584 34.098 ;
        RECT 37.478 34.067 42.538 34.144 ;
        RECT 37.432 34.113 42.492 34.19 ;
        RECT 37.386 34.159 42.446 34.236 ;
        RECT 37.34 34.205 42.4 34.282 ;
        RECT 37.294 34.251 42.354 34.328 ;
        RECT 37.248 34.297 42.308 34.374 ;
        RECT 37.202 34.343 42.262 34.42 ;
        RECT 37.156 34.389 42.216 34.466 ;
        RECT 37.11 34.435 42.17 34.512 ;
        RECT 37.064 34.481 42.124 34.558 ;
        RECT 37.018 34.527 42.078 34.604 ;
        RECT 36.972 34.573 42.032 34.65 ;
        RECT 36.926 34.619 41.986 34.696 ;
        RECT 36.88 34.665 41.94 34.742 ;
        RECT 36.834 34.711 41.894 34.788 ;
        RECT 36.788 34.757 41.848 34.834 ;
        RECT 36.742 34.803 41.802 34.88 ;
        RECT 36.696 34.849 41.756 34.926 ;
        RECT 36.65 34.895 41.71 34.972 ;
        RECT 36.604 34.941 41.664 35.018 ;
        RECT 36.558 34.987 41.618 35.064 ;
        RECT 36.512 35.033 41.572 35.11 ;
        RECT 36.466 35.079 41.526 35.156 ;
        RECT 36.42 35.125 41.48 35.202 ;
        RECT 36.374 35.171 41.434 35.248 ;
        RECT 36.328 35.217 41.388 35.294 ;
        RECT 36.282 35.263 41.342 35.34 ;
        RECT 36.236 35.309 41.296 35.386 ;
        RECT 36.19 35.355 41.25 35.432 ;
        RECT 36.144 35.401 41.204 35.478 ;
        RECT 36.098 35.447 41.158 35.524 ;
        RECT 36.052 35.493 41.112 35.57 ;
        RECT 36.006 35.539 41.066 35.616 ;
        RECT 35.96 35.585 41.02 35.662 ;
        RECT 35.914 35.631 40.974 35.708 ;
        RECT 35.868 35.677 40.928 35.754 ;
        RECT 35.822 35.723 40.882 35.8 ;
        RECT 35.776 35.769 40.836 35.846 ;
        RECT 35.73 35.815 40.79 35.892 ;
        RECT 35.684 35.861 40.744 35.938 ;
        RECT 35.638 35.907 40.698 35.984 ;
        RECT 35.592 35.953 40.652 36.03 ;
        RECT 35.546 35.999 40.606 36.076 ;
        RECT 35.5 36.045 40.56 36.122 ;
        RECT 35.454 36.091 40.514 36.168 ;
        RECT 35.408 36.137 40.468 36.214 ;
        RECT 35.362 36.183 40.422 36.26 ;
        RECT 35.316 36.229 40.376 36.306 ;
        RECT 35.27 36.275 40.33 36.352 ;
        RECT 35.224 36.321 40.284 36.398 ;
        RECT 35.178 36.367 40.238 36.444 ;
        RECT 35.132 36.413 40.192 36.49 ;
        RECT 35.086 36.459 40.146 36.536 ;
        RECT 35.04 36.505 40.1 36.582 ;
        RECT 34.994 36.551 40.054 36.628 ;
        RECT 34.948 36.597 40.008 36.674 ;
        RECT 34.902 36.643 39.962 36.72 ;
        RECT 34.856 36.689 39.916 36.766 ;
        RECT 34.81 36.735 39.87 36.812 ;
        RECT 34.764 36.781 39.824 36.858 ;
        RECT 34.718 36.827 39.778 36.904 ;
        RECT 34.672 36.873 39.732 36.95 ;
        RECT 34.626 36.919 39.686 36.996 ;
        RECT 34.58 36.965 39.64 37.042 ;
        RECT 34.534 37.011 39.594 37.088 ;
        RECT 34.488 37.057 39.548 37.134 ;
        RECT 34.442 37.103 39.502 37.18 ;
        RECT 34.396 37.149 39.456 37.226 ;
        RECT 34.35 37.195 39.41 37.272 ;
        RECT 34.304 37.241 39.364 37.318 ;
        RECT 34.258 37.287 39.318 37.364 ;
        RECT 34.212 37.333 39.272 37.41 ;
        RECT 34.166 37.379 39.226 37.456 ;
        RECT 34.12 37.425 39.18 37.502 ;
        RECT 34.074 37.471 39.134 37.548 ;
        RECT 34.028 37.517 39.088 37.594 ;
        RECT 33.982 37.563 39.042 37.64 ;
        RECT 33.936 37.609 38.996 37.686 ;
        RECT 33.89 37.655 38.95 37.732 ;
        RECT 33.844 37.701 38.904 37.778 ;
        RECT 33.798 37.747 38.858 37.824 ;
        RECT 33.752 37.793 38.812 37.87 ;
        RECT 33.706 37.839 38.766 37.916 ;
        RECT 33.66 37.885 38.72 37.962 ;
        RECT 33.614 37.931 38.674 38.008 ;
        RECT 33.568 37.977 38.628 38.054 ;
        RECT 33.522 38.023 38.582 38.1 ;
        RECT 33.476 38.069 38.536 38.146 ;
        RECT 33.43 38.115 38.49 38.192 ;
        RECT 33.384 38.161 38.444 38.238 ;
        RECT 33.338 38.207 38.398 38.284 ;
        RECT 33.292 38.253 38.352 38.33 ;
        RECT 33.246 38.299 38.306 38.376 ;
        RECT 33.2 38.345 38.26 38.422 ;
        RECT 33.154 38.391 38.214 38.468 ;
        RECT 33.108 38.437 38.168 38.514 ;
        RECT 33.062 38.483 38.122 38.56 ;
        RECT 33.016 38.529 38.076 38.606 ;
        RECT 32.97 38.575 38.03 38.652 ;
        RECT 32.924 38.621 37.984 38.698 ;
        RECT 32.878 38.667 37.938 38.744 ;
        RECT 32.832 38.713 37.892 38.79 ;
        RECT 32.786 38.759 37.846 38.836 ;
        RECT 32.74 38.805 37.8 38.882 ;
        RECT 32.694 38.851 37.754 38.928 ;
        RECT 32.648 38.897 37.708 38.974 ;
        RECT 32.602 38.943 37.662 39.02 ;
        RECT 32.556 38.989 37.616 39.066 ;
        RECT 32.51 39.035 37.57 39.112 ;
        RECT 32.464 39.081 37.524 39.158 ;
        RECT 32.418 39.127 37.478 39.204 ;
        RECT 32.372 39.173 37.432 39.25 ;
        RECT 32.326 39.219 37.386 39.296 ;
        RECT 32.28 39.265 37.34 39.342 ;
        RECT 32.234 39.311 37.294 39.388 ;
        RECT 32.188 39.357 37.248 39.434 ;
        RECT 32.142 39.403 37.202 39.48 ;
        RECT 32.096 39.449 37.156 39.526 ;
        RECT 32.05 39.495 37.11 39.572 ;
        RECT 32.004 39.541 37.064 39.618 ;
        RECT 31.958 39.587 37.018 39.664 ;
        RECT 31.912 39.633 36.972 39.71 ;
        RECT 31.866 39.679 36.926 39.756 ;
        RECT 31.82 39.725 36.88 39.802 ;
        RECT 31.774 39.771 36.834 39.848 ;
        RECT 31.728 39.817 36.788 39.894 ;
        RECT 31.682 39.863 36.742 39.94 ;
        RECT 31.636 39.909 36.696 39.986 ;
        RECT 31.59 39.955 36.65 40.032 ;
        RECT 31.544 40.001 36.604 40.078 ;
        RECT 31.498 40.047 36.558 40.124 ;
        RECT 31.452 40.093 36.512 40.17 ;
        RECT 31.406 40.139 36.466 40.216 ;
        RECT 31.36 40.185 36.42 40.262 ;
        RECT 31.314 40.231 36.374 40.308 ;
        RECT 31.268 40.277 36.328 40.354 ;
        RECT 31.222 40.323 36.282 40.4 ;
        RECT 31.176 40.369 36.236 40.446 ;
        RECT 31.13 40.415 36.19 40.492 ;
        RECT 31.084 40.461 36.144 40.538 ;
        RECT 31.038 40.507 36.098 40.584 ;
        RECT 30.992 40.553 36.052 40.63 ;
        RECT 30.946 40.599 36.006 40.676 ;
        RECT 30.9 40.645 35.96 40.722 ;
        RECT 30.854 40.691 35.914 40.768 ;
        RECT 30.808 40.737 35.868 40.814 ;
        RECT 30.762 40.783 35.822 40.86 ;
        RECT 30.716 40.829 35.776 40.906 ;
        RECT 30.67 40.875 35.73 40.952 ;
        RECT 30.624 40.921 35.684 40.998 ;
        RECT 30.578 40.967 35.638 41.044 ;
        RECT 30.532 41.013 35.592 41.09 ;
        RECT 30.486 41.059 35.546 41.136 ;
        RECT 30.44 41.105 35.5 41.182 ;
        RECT 30.394 41.151 35.454 41.228 ;
        RECT 30.348 41.197 35.408 41.274 ;
        RECT 30.302 41.243 35.362 41.32 ;
        RECT 30.256 41.289 35.316 41.366 ;
        RECT 30.21 41.335 35.27 41.412 ;
        RECT 30.164 41.381 35.224 41.458 ;
        RECT 30.118 41.427 35.178 41.504 ;
        RECT 30.072 41.473 35.132 41.55 ;
        RECT 30.026 41.519 35.086 41.596 ;
        RECT 29.98 41.565 35.04 41.642 ;
        RECT 29.934 41.611 34.994 41.688 ;
        RECT 29.888 41.657 34.948 41.734 ;
        RECT 29.842 41.703 34.902 41.78 ;
        RECT 29.796 41.749 34.856 41.826 ;
        RECT 29.75 41.795 34.81 41.872 ;
        RECT 29.704 41.841 34.764 41.918 ;
        RECT 29.658 41.887 34.718 41.964 ;
        RECT 29.612 41.933 34.672 42.01 ;
        RECT 29.566 41.979 34.626 42.056 ;
        RECT 29.52 42.025 34.58 42.102 ;
        RECT 29.474 42.071 34.534 42.148 ;
        RECT 29.428 42.117 34.488 42.194 ;
        RECT 29.382 42.163 34.442 42.24 ;
        RECT 29.336 42.209 34.396 42.286 ;
        RECT 29.29 42.255 34.35 42.332 ;
        RECT 29.244 42.301 34.304 42.378 ;
        RECT 29.198 42.347 34.258 42.424 ;
        RECT 29.152 42.393 34.212 42.47 ;
        RECT 29.106 42.439 34.166 42.516 ;
        RECT 29.06 42.485 34.12 42.562 ;
        RECT 29.014 42.531 34.074 42.608 ;
        RECT 28.968 42.577 34.028 42.654 ;
        RECT 28.922 42.623 33.982 42.7 ;
        RECT 28.876 42.669 33.936 42.746 ;
        RECT 28.83 42.715 33.89 42.792 ;
        RECT 28.784 42.761 33.844 42.838 ;
        RECT 28.738 42.807 33.798 42.884 ;
        RECT 28.692 42.853 33.752 42.93 ;
        RECT 28.646 42.899 33.706 42.976 ;
        RECT 28.6 42.945 33.66 43.022 ;
        RECT 28.554 42.991 33.614 43.068 ;
        RECT 28.508 43.037 33.568 43.114 ;
        RECT 28.462 43.083 33.522 43.16 ;
        RECT 28.416 43.129 33.476 43.206 ;
        RECT 28.37 43.175 33.43 43.252 ;
        RECT 28.324 43.221 33.384 43.298 ;
        RECT 28.278 43.267 33.338 43.344 ;
        RECT 28.232 43.313 33.292 43.39 ;
        RECT 28.186 43.359 33.246 43.436 ;
        RECT 28.14 43.405 33.2 43.482 ;
        RECT 28.094 43.451 33.154 43.528 ;
        RECT 28.048 43.497 33.108 43.574 ;
        RECT 28.002 43.543 33.062 43.62 ;
        RECT 27.956 43.589 33.016 43.666 ;
        RECT 27.91 43.635 32.97 43.712 ;
        RECT 27.864 43.681 32.924 43.758 ;
        RECT 27.818 43.727 32.878 43.804 ;
        RECT 27.772 43.773 32.832 43.85 ;
        RECT 27.726 43.819 32.786 43.896 ;
        RECT 27.68 43.865 32.74 43.942 ;
        RECT 27.634 43.911 32.694 43.988 ;
        RECT 27.588 43.957 32.648 44.034 ;
        RECT 27.542 44.003 32.602 44.08 ;
        RECT 27.496 44.049 32.556 44.126 ;
        RECT 27.45 44.095 32.51 44.172 ;
        RECT 27.404 44.141 32.464 44.218 ;
        RECT 27.358 44.187 32.418 44.264 ;
        RECT 27.312 44.233 32.372 44.31 ;
        RECT 27.266 44.279 32.326 44.356 ;
        RECT 27.22 44.325 32.28 44.402 ;
        RECT 27.174 44.371 32.234 44.448 ;
        RECT 27.128 44.417 32.188 44.494 ;
        RECT 27.082 44.463 32.142 44.54 ;
        RECT 27.036 44.509 32.096 44.586 ;
        RECT 26.99 44.555 32.05 44.632 ;
        RECT 26.944 44.601 32.004 44.678 ;
        RECT 26.898 44.647 31.958 44.724 ;
        RECT 26.852 44.693 31.912 44.77 ;
        RECT 26.806 44.739 31.866 44.816 ;
        RECT 26.76 44.785 31.82 44.862 ;
        RECT 26.714 44.831 31.774 44.908 ;
        RECT 26.668 44.877 31.728 44.954 ;
        RECT 26.622 44.923 31.682 45 ;
        RECT 26.576 44.969 31.636 45.046 ;
        RECT 26.53 45.015 31.59 45.092 ;
        RECT 26.484 45.061 31.544 45.138 ;
        RECT 26.438 45.107 31.498 45.184 ;
        RECT 26.392 45.153 31.452 45.23 ;
        RECT 26.346 45.199 31.406 45.276 ;
        RECT 26.3 45.245 31.36 45.322 ;
        RECT 26.254 45.291 31.314 45.368 ;
        RECT 26.208 45.337 31.268 45.414 ;
        RECT 26.162 45.383 31.222 45.46 ;
        RECT 26.116 45.429 31.176 45.506 ;
        RECT 26.07 45.475 31.13 45.552 ;
        RECT 26.024 45.521 31.084 45.598 ;
        RECT 25.978 45.567 31.038 45.644 ;
        RECT 25.932 45.613 30.992 45.69 ;
        RECT 25.886 45.659 30.946 45.736 ;
        RECT 25.84 45.705 30.9 45.782 ;
        RECT 25.794 45.751 30.854 45.828 ;
        RECT 25.748 45.797 30.808 45.874 ;
        RECT 25.702 45.843 30.762 45.92 ;
        RECT 25.656 45.889 30.716 45.966 ;
        RECT 25.61 45.935 30.67 46.012 ;
        RECT 25.564 45.981 30.624 46.058 ;
        RECT 25.518 46.027 30.578 46.104 ;
        RECT 25.472 46.073 30.532 46.15 ;
        RECT 25.426 46.119 30.486 46.196 ;
        RECT 25.38 46.165 30.44 46.242 ;
        RECT 25.334 46.211 30.394 46.288 ;
        RECT 25.288 46.257 30.348 46.334 ;
        RECT 25.242 46.303 30.302 46.38 ;
        RECT 25.196 46.349 30.256 46.426 ;
        RECT 25.15 46.395 30.21 46.472 ;
        RECT 25.104 46.441 30.164 46.518 ;
        RECT 25.058 46.487 30.118 46.564 ;
        RECT 25.012 46.533 30.072 46.61 ;
        RECT 24.966 46.579 30.026 46.656 ;
        RECT 24.92 46.625 29.98 46.702 ;
        RECT 24.874 46.671 29.934 46.748 ;
        RECT 24.828 46.717 29.888 46.794 ;
        RECT 24.782 46.763 29.842 46.84 ;
        RECT 24.736 46.809 29.796 46.886 ;
        RECT 24.69 46.855 29.75 46.932 ;
        RECT 24.644 46.901 29.704 46.978 ;
        RECT 24.598 46.947 29.658 47.024 ;
        RECT 24.552 46.993 29.612 47.07 ;
        RECT 24.506 47.039 29.566 47.116 ;
        RECT 24.46 47.085 29.52 47.162 ;
        RECT 24.414 47.131 29.474 47.208 ;
        RECT 24.368 47.177 29.428 47.254 ;
        RECT 24.322 47.223 29.382 47.3 ;
        RECT 24.276 47.269 29.336 47.346 ;
        RECT 24.23 47.315 29.29 47.392 ;
        RECT 24.184 47.361 29.244 47.438 ;
        RECT 24.138 47.407 29.198 47.484 ;
        RECT 24.092 47.453 29.152 47.53 ;
        RECT 24.046 47.499 29.106 47.576 ;
        RECT 24 47.545 29.06 47.622 ;
        RECT 23.954 47.591 29.014 47.668 ;
        RECT 23.908 47.637 28.968 47.714 ;
        RECT 23.862 47.683 28.922 47.76 ;
        RECT 23.816 47.729 28.876 47.806 ;
        RECT 23.77 47.775 28.83 47.852 ;
        RECT 23.724 47.821 28.784 47.898 ;
        RECT 23.678 47.867 28.738 47.944 ;
        RECT 23.632 47.913 28.692 47.99 ;
        RECT 23.586 47.959 28.646 48.036 ;
        RECT 23.54 48.005 28.6 48.082 ;
        RECT 23.494 48.051 28.554 48.128 ;
        RECT 23.448 48.097 28.508 48.174 ;
        RECT 23.402 48.143 28.462 48.22 ;
        RECT 23.356 48.189 28.416 48.266 ;
        RECT 23.31 48.235 28.37 48.312 ;
        RECT 23.264 48.281 28.324 48.358 ;
        RECT 23.218 48.327 28.278 48.404 ;
        RECT 23.172 48.373 28.232 48.45 ;
        RECT 23.126 48.419 28.186 48.496 ;
        RECT 23.08 48.465 28.14 48.542 ;
        RECT 23.034 48.511 28.094 48.588 ;
        RECT 22.988 48.557 28.048 48.634 ;
        RECT 22.942 48.603 28.002 48.68 ;
        RECT 22.896 48.649 27.956 48.726 ;
        RECT 22.85 48.695 27.91 48.772 ;
        RECT 22.804 48.741 27.864 48.818 ;
        RECT 22.758 48.787 27.818 48.864 ;
        RECT 22.712 48.833 27.772 48.91 ;
        RECT 22.666 48.879 27.726 48.956 ;
        RECT 22.62 48.925 27.68 49.002 ;
        RECT 22.574 48.971 27.634 49.048 ;
        RECT 22.528 49.017 27.588 49.094 ;
        RECT 22.482 49.063 27.542 49.14 ;
        RECT 22.436 49.109 27.496 49.186 ;
        RECT 22.39 49.155 27.45 49.232 ;
        RECT 22.344 49.201 27.404 49.278 ;
        RECT 22.298 49.247 27.358 49.324 ;
        RECT 22.252 49.293 27.312 49.37 ;
        RECT 22.206 49.339 27.266 49.416 ;
        RECT 22.16 49.385 27.22 49.462 ;
        RECT 22.114 49.431 27.174 49.508 ;
        RECT 22.068 49.477 27.128 49.554 ;
        RECT 22.022 49.523 27.082 49.6 ;
        RECT 21.976 49.569 27.036 49.646 ;
        RECT 21.93 49.615 26.99 49.692 ;
        RECT 21.884 49.661 26.944 49.738 ;
        RECT 21.838 49.707 26.898 49.784 ;
        RECT 21.792 49.753 26.852 49.83 ;
        RECT 21.746 49.799 26.806 49.876 ;
        RECT 21.7 49.845 26.76 49.922 ;
        RECT 21.654 49.891 26.714 49.968 ;
        RECT 21.608 49.937 26.668 50.014 ;
        RECT 21.562 49.983 26.622 50.06 ;
        RECT 21.516 50.029 26.576 50.106 ;
        RECT 21.47 50.075 26.53 50.152 ;
        RECT 21.424 50.121 26.484 50.198 ;
        RECT 21.378 50.167 26.438 50.244 ;
        RECT 21.332 50.213 26.392 50.29 ;
        RECT 21.286 50.259 26.346 50.336 ;
        RECT 21.24 50.305 26.3 50.382 ;
        RECT 21.194 50.351 26.254 50.428 ;
        RECT 21.148 50.397 26.208 50.474 ;
        RECT 21.102 50.443 26.162 50.52 ;
        RECT 21.056 50.489 26.116 50.566 ;
        RECT 21.01 50.535 26.07 50.612 ;
        RECT 20.964 50.581 26.024 50.658 ;
        RECT 20.918 50.627 25.978 50.704 ;
        RECT 20.872 50.673 25.932 50.75 ;
        RECT 20.826 50.719 25.886 50.796 ;
        RECT 20.78 50.765 25.84 50.842 ;
        RECT 20.734 50.811 25.794 50.888 ;
        RECT 20.688 50.857 25.748 50.934 ;
        RECT 20.642 50.903 25.702 50.98 ;
        RECT 20.596 50.949 25.656 51.026 ;
        RECT 20.55 50.995 25.61 51.072 ;
        RECT 20.504 51.041 25.564 51.118 ;
        RECT 20.458 51.087 25.518 51.164 ;
        RECT 20.412 51.133 25.472 51.21 ;
        RECT 20.366 51.179 25.426 51.256 ;
        RECT 20.32 51.225 25.38 51.302 ;
        RECT 20.274 51.271 25.334 51.348 ;
        RECT 20.228 51.317 25.288 51.394 ;
        RECT 20.182 51.363 25.242 51.44 ;
        RECT 20.136 51.409 25.196 51.486 ;
        RECT 20.09 51.455 25.15 51.532 ;
        RECT 20.044 51.501 25.104 51.578 ;
        RECT 19.998 51.547 25.058 51.624 ;
        RECT 19.952 51.593 25.012 51.67 ;
        RECT 19.906 51.639 24.966 51.716 ;
        RECT 19.86 51.685 24.92 51.762 ;
        RECT 19.814 51.731 24.874 51.808 ;
        RECT 19.768 51.777 24.828 51.854 ;
        RECT 19.722 51.823 24.782 51.9 ;
        RECT 19.676 51.869 24.736 51.946 ;
        RECT 19.63 51.915 24.69 51.992 ;
        RECT 19.584 51.961 24.644 52.038 ;
        RECT 19.538 52.007 24.598 52.084 ;
        RECT 19.492 52.053 24.552 52.13 ;
        RECT 19.446 52.099 24.506 52.176 ;
        RECT 19.4 52.145 24.46 52.222 ;
        RECT 19.354 52.191 24.414 52.268 ;
        RECT 19.308 52.237 24.368 52.314 ;
        RECT 19.262 52.283 24.322 52.36 ;
        RECT 19.216 52.329 24.276 52.406 ;
        RECT 19.17 52.375 24.23 52.452 ;
        RECT 19.124 52.421 24.184 52.498 ;
        RECT 19.078 52.467 24.138 52.544 ;
        RECT 19.032 52.513 24.092 52.59 ;
        RECT 18.986 52.559 24.046 52.636 ;
        RECT 18.94 52.605 24 52.682 ;
        RECT 18.894 52.651 23.954 52.728 ;
        RECT 18.848 52.697 23.908 52.774 ;
        RECT 18.802 52.743 23.862 52.82 ;
        RECT 18.756 52.789 23.816 52.866 ;
        RECT 18.71 52.835 23.77 52.912 ;
        RECT 18.664 52.881 23.724 52.958 ;
        RECT 18.618 52.927 23.678 53.004 ;
        RECT 18.572 52.973 23.632 53.05 ;
    END
    PORT
      LAYER IB ;
        RECT 68.154 49.95 80 53.55 ;
        RECT 64.544 53.537 69.645 53.56 ;
        RECT 63.118 54.963 68.2 55.018 ;
        RECT 68.132 49.961 68.154 55.052 ;
        RECT 63.072 55.009 68.132 55.086 ;
        RECT 63.164 54.917 68.246 54.972 ;
        RECT 68.086 49.995 68.132 55.086 ;
        RECT 63.026 55.055 68.086 55.132 ;
        RECT 63.21 54.871 68.292 54.926 ;
        RECT 68.04 50.041 68.086 55.132 ;
        RECT 62.98 55.101 68.04 55.178 ;
        RECT 63.256 54.825 68.338 54.88 ;
        RECT 67.994 50.087 68.04 55.178 ;
        RECT 62.934 55.147 67.994 55.224 ;
        RECT 63.302 54.779 68.384 54.834 ;
        RECT 67.948 50.133 67.994 55.224 ;
        RECT 62.888 55.193 67.948 55.27 ;
        RECT 63.348 54.733 68.43 54.788 ;
        RECT 67.902 50.179 67.948 55.27 ;
        RECT 62.842 55.239 67.902 55.316 ;
        RECT 63.394 54.687 68.476 54.742 ;
        RECT 67.856 50.225 67.902 55.316 ;
        RECT 62.796 55.285 67.856 55.362 ;
        RECT 63.44 54.641 68.522 54.696 ;
        RECT 67.81 50.271 67.856 55.362 ;
        RECT 62.75 55.331 67.81 55.408 ;
        RECT 63.486 54.595 68.568 54.65 ;
        RECT 67.764 50.317 67.81 55.408 ;
        RECT 62.704 55.377 67.764 55.454 ;
        RECT 63.532 54.549 68.614 54.604 ;
        RECT 67.718 50.363 67.764 55.454 ;
        RECT 62.658 55.423 67.718 55.5 ;
        RECT 63.578 54.503 68.66 54.558 ;
        RECT 67.672 50.409 67.718 55.5 ;
        RECT 62.612 55.469 67.672 55.546 ;
        RECT 63.624 54.457 68.706 54.512 ;
        RECT 67.626 50.455 67.672 55.546 ;
        RECT 62.566 55.515 67.626 55.592 ;
        RECT 63.67 54.411 68.752 54.466 ;
        RECT 67.58 50.501 67.626 55.592 ;
        RECT 62.52 55.561 67.58 55.638 ;
        RECT 63.716 54.365 68.798 54.42 ;
        RECT 67.534 50.547 67.58 55.638 ;
        RECT 62.474 55.607 67.534 55.684 ;
        RECT 63.762 54.319 68.844 54.374 ;
        RECT 67.488 50.593 67.534 55.684 ;
        RECT 62.428 55.653 67.488 55.73 ;
        RECT 63.808 54.273 68.89 54.328 ;
        RECT 67.442 50.639 67.488 55.73 ;
        RECT 62.382 55.699 67.442 55.776 ;
        RECT 63.854 54.227 68.936 54.282 ;
        RECT 67.396 50.685 67.442 55.776 ;
        RECT 62.336 55.745 67.396 55.822 ;
        RECT 63.9 54.181 68.982 54.236 ;
        RECT 67.35 50.731 67.396 55.822 ;
        RECT 62.29 55.791 67.35 55.868 ;
        RECT 63.946 54.135 69.028 54.19 ;
        RECT 67.304 50.777 67.35 55.868 ;
        RECT 62.244 55.837 67.304 55.914 ;
        RECT 63.992 54.089 69.074 54.144 ;
        RECT 67.258 50.823 67.304 55.914 ;
        RECT 62.198 55.883 67.258 55.96 ;
        RECT 64.038 54.043 69.12 54.098 ;
        RECT 67.212 50.869 67.258 55.96 ;
        RECT 62.152 55.929 67.212 56.006 ;
        RECT 64.084 53.997 69.166 54.052 ;
        RECT 67.166 50.915 67.212 56.006 ;
        RECT 62.106 55.975 67.166 56.052 ;
        RECT 64.13 53.951 69.212 54.006 ;
        RECT 67.12 50.961 67.166 56.052 ;
        RECT 62.06 56.021 67.12 56.098 ;
        RECT 64.176 53.905 69.258 53.96 ;
        RECT 67.074 51.007 67.12 56.098 ;
        RECT 62.014 56.067 67.074 56.144 ;
        RECT 64.222 53.859 69.304 53.914 ;
        RECT 67.028 51.053 67.074 56.144 ;
        RECT 61.968 56.113 67.028 56.19 ;
        RECT 64.268 53.813 69.35 53.868 ;
        RECT 66.982 51.099 67.028 56.19 ;
        RECT 61.922 56.159 66.982 56.236 ;
        RECT 64.314 53.767 69.396 53.822 ;
        RECT 66.936 51.145 66.982 56.236 ;
        RECT 61.876 56.205 66.936 56.282 ;
        RECT 64.36 53.721 69.442 53.776 ;
        RECT 66.89 51.191 66.936 56.282 ;
        RECT 61.83 56.251 66.89 56.328 ;
        RECT 64.406 53.675 69.488 53.73 ;
        RECT 66.844 51.237 66.89 56.328 ;
        RECT 61.784 56.297 66.844 56.374 ;
        RECT 64.452 53.629 69.534 53.684 ;
        RECT 66.798 51.283 66.844 56.374 ;
        RECT 61.738 56.343 66.798 56.42 ;
        RECT 64.498 53.583 69.58 53.638 ;
        RECT 66.752 51.329 66.798 56.42 ;
        RECT 61.692 56.389 66.752 56.466 ;
        RECT 64.544 53.537 69.626 53.592 ;
        RECT 66.706 51.375 66.752 56.466 ;
        RECT 61.646 56.435 66.706 56.512 ;
        RECT 64.59 53.491 80 53.55 ;
        RECT 66.66 51.421 66.706 56.512 ;
        RECT 61.6 56.481 66.66 56.558 ;
        RECT 64.636 53.445 80 53.55 ;
        RECT 66.614 51.467 66.66 56.558 ;
        RECT 61.554 56.527 66.614 56.604 ;
        RECT 64.682 53.399 80 53.55 ;
        RECT 66.568 51.513 66.614 56.604 ;
        RECT 61.508 56.573 66.568 56.65 ;
        RECT 64.728 53.353 80 53.55 ;
        RECT 66.522 51.559 66.568 56.65 ;
        RECT 61.462 56.619 66.522 56.696 ;
        RECT 64.774 53.307 80 53.55 ;
        RECT 66.476 51.605 66.522 56.696 ;
        RECT 61.416 56.665 66.476 56.742 ;
        RECT 64.82 53.261 80 53.55 ;
        RECT 66.43 51.651 66.476 56.742 ;
        RECT 61.37 56.711 66.43 56.788 ;
        RECT 64.866 53.215 80 53.55 ;
        RECT 66.384 51.697 66.43 56.788 ;
        RECT 61.324 56.757 66.384 56.834 ;
        RECT 64.912 53.169 80 53.55 ;
        RECT 66.338 51.743 66.384 56.834 ;
        RECT 61.278 56.803 66.338 56.88 ;
        RECT 64.958 53.123 80 53.55 ;
        RECT 66.292 51.789 66.338 56.88 ;
        RECT 61.232 56.849 66.292 56.926 ;
        RECT 65.004 53.077 80 53.55 ;
        RECT 66.246 51.835 66.292 56.926 ;
        RECT 61.186 56.895 66.246 56.972 ;
        RECT 65.05 53.031 80 53.55 ;
        RECT 66.2 51.881 66.246 56.972 ;
        RECT 61.14 56.941 66.2 57.018 ;
        RECT 65.096 52.985 80 53.55 ;
        RECT 66.154 51.927 66.2 57.018 ;
        RECT 61.094 56.987 66.154 57.064 ;
        RECT 65.142 52.939 80 53.55 ;
        RECT 66.108 51.973 66.154 57.064 ;
        RECT 61.048 57.033 66.108 57.11 ;
        RECT 65.188 52.893 80 53.55 ;
        RECT 66.062 52.019 66.108 57.11 ;
        RECT 61.002 57.079 66.062 57.156 ;
        RECT 65.234 52.847 80 53.55 ;
        RECT 66.016 52.065 66.062 57.156 ;
        RECT 60.956 57.125 66.016 57.202 ;
        RECT 65.28 52.801 80 53.55 ;
        RECT 65.97 52.111 66.016 57.202 ;
        RECT 60.91 57.171 65.97 57.248 ;
        RECT 65.326 52.755 80 53.55 ;
        RECT 65.924 52.157 65.97 57.248 ;
        RECT 60.864 57.217 65.924 57.294 ;
        RECT 65.372 52.709 80 53.55 ;
        RECT 65.878 52.203 65.924 57.294 ;
        RECT 60.818 57.263 65.878 57.34 ;
        RECT 65.418 52.663 80 53.55 ;
        RECT 65.832 52.249 65.878 57.34 ;
        RECT 60.772 57.309 65.832 57.386 ;
        RECT 65.464 52.617 80 53.55 ;
        RECT 65.786 52.295 65.832 57.386 ;
        RECT 60.726 57.355 65.786 57.432 ;
        RECT 65.51 52.571 80 53.55 ;
        RECT 65.74 52.341 65.786 57.432 ;
        RECT 60.68 57.401 65.74 57.478 ;
        RECT 65.556 52.525 80 53.55 ;
        RECT 65.694 52.387 65.74 57.478 ;
        RECT 60.634 57.447 65.694 57.524 ;
        RECT 65.602 52.479 80 53.55 ;
        RECT 65.648 52.433 65.694 57.524 ;
        RECT 60.588 57.493 65.648 57.57 ;
        RECT 60.542 57.539 65.602 57.616 ;
        RECT 60.496 57.585 65.556 57.662 ;
        RECT 60.45 57.631 65.51 57.708 ;
        RECT 60.404 57.677 65.464 57.754 ;
        RECT 60.358 57.723 65.418 57.8 ;
        RECT 60.312 57.769 65.372 57.846 ;
        RECT 60.266 57.815 65.326 57.892 ;
        RECT 60.22 57.861 65.28 57.938 ;
        RECT 60.174 57.907 65.234 57.984 ;
        RECT 60.128 57.953 65.188 58.03 ;
        RECT 60.082 57.999 65.142 58.076 ;
        RECT 60.036 58.045 65.096 58.122 ;
        RECT 59.99 58.091 65.05 58.168 ;
        RECT 59.944 58.137 65.004 58.214 ;
        RECT 59.898 58.183 64.958 58.26 ;
        RECT 59.852 58.229 64.912 58.306 ;
        RECT 59.806 58.275 64.866 58.352 ;
        RECT 59.76 58.321 64.82 58.398 ;
        RECT 59.714 58.367 64.774 58.444 ;
        RECT 59.668 58.413 64.728 58.49 ;
        RECT 59.622 58.459 64.682 58.536 ;
        RECT 59.576 58.505 64.636 58.582 ;
        RECT 59.53 58.551 64.59 58.628 ;
        RECT 59.484 58.597 64.544 58.674 ;
        RECT 59.438 58.643 64.498 58.72 ;
        RECT 59.392 58.689 64.452 58.766 ;
        RECT 59.346 58.735 64.406 58.812 ;
        RECT 59.3 58.781 64.36 58.858 ;
        RECT 59.254 58.827 64.314 58.904 ;
        RECT 59.208 58.873 64.268 58.95 ;
        RECT 59.162 58.919 64.222 58.996 ;
        RECT 59.116 58.965 64.176 59.042 ;
        RECT 59.07 59.011 64.13 59.088 ;
        RECT 59.024 59.057 64.084 59.134 ;
        RECT 58.978 59.103 64.038 59.18 ;
        RECT 58.932 59.149 63.992 59.226 ;
        RECT 58.886 59.195 63.946 59.272 ;
        RECT 58.84 59.241 63.9 59.318 ;
        RECT 58.794 59.287 63.854 59.364 ;
        RECT 58.748 59.333 63.808 59.41 ;
        RECT 58.702 59.379 63.762 59.456 ;
        RECT 58.656 59.425 63.716 59.502 ;
        RECT 58.61 59.471 63.67 59.548 ;
        RECT 58.564 59.517 63.624 59.594 ;
        RECT 58.518 59.563 63.578 59.64 ;
        RECT 58.472 59.609 63.532 59.686 ;
        RECT 58.426 59.655 63.486 59.732 ;
        RECT 58.38 59.701 63.44 59.778 ;
        RECT 58.334 59.747 63.394 59.824 ;
        RECT 58.288 59.793 63.348 59.87 ;
        RECT 58.242 59.839 63.302 59.916 ;
        RECT 58.196 59.885 63.256 59.962 ;
        RECT 58.15 59.931 63.21 60.008 ;
        RECT 58.104 59.977 63.164 60.054 ;
        RECT 58.058 60.023 63.118 60.1 ;
        RECT 58.012 60.069 63.072 60.146 ;
        RECT 57.966 60.115 63.026 60.192 ;
        RECT 57.92 60.161 62.98 60.238 ;
        RECT 57.874 60.207 62.934 60.284 ;
        RECT 57.828 60.253 62.888 60.33 ;
        RECT 57.782 60.299 62.842 60.376 ;
        RECT 57.736 60.345 62.796 60.422 ;
        RECT 57.69 60.391 62.75 60.468 ;
        RECT 57.644 60.437 62.704 60.514 ;
        RECT 57.598 60.483 62.658 60.56 ;
        RECT 57.552 60.529 62.612 60.606 ;
        RECT 57.506 60.575 62.566 60.652 ;
        RECT 57.46 60.621 62.52 60.698 ;
        RECT 57.414 60.667 62.474 60.744 ;
        RECT 57.368 60.713 62.428 60.79 ;
        RECT 57.322 60.759 62.382 60.836 ;
        RECT 57.276 60.805 62.336 60.882 ;
        RECT 57.23 60.851 62.29 60.928 ;
        RECT 57.184 60.897 62.244 60.974 ;
        RECT 57.138 60.943 62.198 61.02 ;
        RECT 57.092 60.989 62.152 61.066 ;
        RECT 57.046 61.035 62.106 61.112 ;
        RECT 57 61.081 62.06 61.158 ;
        RECT 56.954 61.127 62.014 61.204 ;
        RECT 56.908 61.173 61.968 61.25 ;
        RECT 56.862 61.219 61.922 61.296 ;
        RECT 56.816 61.265 61.876 61.342 ;
        RECT 56.77 61.311 61.83 61.388 ;
        RECT 56.724 61.357 61.784 61.434 ;
        RECT 56.678 61.403 61.738 61.48 ;
        RECT 56.632 61.449 61.692 61.526 ;
        RECT 56.586 61.495 61.646 61.572 ;
        RECT 56.54 61.541 61.6 61.618 ;
        RECT 56.494 61.587 61.554 61.664 ;
        RECT 56.448 61.633 61.508 61.71 ;
        RECT 56.402 61.679 61.462 61.756 ;
        RECT 56.356 61.725 61.416 61.802 ;
        RECT 56.31 61.771 61.37 61.848 ;
        RECT 56.264 61.817 61.324 61.894 ;
        RECT 56.218 61.863 61.278 61.94 ;
        RECT 56.172 61.909 61.232 61.986 ;
        RECT 56.126 61.955 61.186 62.032 ;
        RECT 56.08 62.001 61.14 62.078 ;
        RECT 56.034 62.047 61.094 62.124 ;
        RECT 55.988 62.093 61.048 62.17 ;
        RECT 55.942 62.139 61.002 62.216 ;
        RECT 55.896 62.185 60.956 62.262 ;
        RECT 55.85 62.231 60.91 62.308 ;
        RECT 55.804 62.277 60.864 62.354 ;
        RECT 55.758 62.323 60.818 62.4 ;
        RECT 55.712 62.369 60.772 62.446 ;
        RECT 55.666 62.415 60.726 62.492 ;
        RECT 55.62 62.461 60.68 62.538 ;
        RECT 55.574 62.507 60.634 62.584 ;
        RECT 55.528 62.553 60.588 62.63 ;
        RECT 55.482 62.599 60.542 62.676 ;
        RECT 55.436 62.645 60.496 62.722 ;
        RECT 55.39 62.691 60.45 62.768 ;
        RECT 55.344 62.737 60.404 62.814 ;
        RECT 55.298 62.783 60.358 62.86 ;
        RECT 55.252 62.829 60.312 62.906 ;
        RECT 55.206 62.875 60.266 62.952 ;
        RECT 55.16 62.921 60.22 62.998 ;
        RECT 55.114 62.967 60.174 63.044 ;
        RECT 55.068 63.013 60.128 63.09 ;
        RECT 55.022 63.059 60.082 63.136 ;
        RECT 54.976 63.105 60.036 63.182 ;
        RECT 54.93 63.151 59.99 63.228 ;
        RECT 54.884 63.197 59.944 63.274 ;
        RECT 54.838 63.243 59.898 63.32 ;
        RECT 54.792 63.289 59.852 63.366 ;
        RECT 54.746 63.335 59.806 63.412 ;
        RECT 54.7 63.381 59.76 63.458 ;
        RECT 54.654 63.427 59.714 63.504 ;
        RECT 54.608 63.473 59.668 63.55 ;
        RECT 54.562 63.519 59.622 63.596 ;
        RECT 54.516 63.565 59.576 63.642 ;
        RECT 54.47 63.611 59.53 63.688 ;
        RECT 54.424 63.657 59.484 63.734 ;
        RECT 54.378 63.703 59.438 63.78 ;
        RECT 54.332 63.749 59.392 63.826 ;
        RECT 54.286 63.795 59.346 63.872 ;
        RECT 54.24 63.841 59.3 63.918 ;
        RECT 54.194 63.887 59.254 63.964 ;
        RECT 54.148 63.933 59.208 64.01 ;
        RECT 54.102 63.979 59.162 64.056 ;
        RECT 54.056 64.025 59.116 64.102 ;
        RECT 54.01 64.071 59.07 64.148 ;
        RECT 53.964 64.117 59.024 64.194 ;
        RECT 53.918 64.163 58.978 64.24 ;
        RECT 53.872 64.209 58.932 64.286 ;
        RECT 53.826 64.255 58.886 64.332 ;
        RECT 53.78 64.301 58.84 64.378 ;
        RECT 53.734 64.347 58.794 64.424 ;
        RECT 53.688 64.393 58.748 64.47 ;
        RECT 53.642 64.439 58.702 64.516 ;
        RECT 53.55 64.531 58.656 64.562 ;
        RECT 53.596 64.485 58.656 64.562 ;
        RECT 53.538 64.56 58.61 64.608 ;
        RECT 53.492 64.589 58.564 64.654 ;
        RECT 53.446 64.635 58.518 64.7 ;
        RECT 53.4 64.681 58.472 64.746 ;
        RECT 53.354 64.727 58.426 64.792 ;
        RECT 53.308 64.773 58.38 64.838 ;
        RECT 53.262 64.819 58.334 64.884 ;
        RECT 53.216 64.865 58.288 64.93 ;
        RECT 53.17 64.911 58.242 64.976 ;
        RECT 53.124 64.957 58.196 65.022 ;
        RECT 53.078 65.003 58.15 65.068 ;
        RECT 53.032 65.049 58.104 65.114 ;
        RECT 52.986 65.095 58.058 65.16 ;
        RECT 52.94 65.141 58.012 65.206 ;
        RECT 52.894 65.187 57.966 65.252 ;
        RECT 52.848 65.233 57.92 65.298 ;
        RECT 52.802 65.279 57.874 65.344 ;
        RECT 52.756 65.325 57.828 65.39 ;
        RECT 52.71 65.371 57.782 65.436 ;
        RECT 52.664 65.417 57.736 65.482 ;
        RECT 52.618 65.463 57.69 65.528 ;
        RECT 52.572 65.509 57.644 65.574 ;
        RECT 52.526 65.555 57.598 65.62 ;
        RECT 52.48 65.601 57.552 65.666 ;
        RECT 52.434 65.647 57.506 65.712 ;
        RECT 52.388 65.693 57.46 65.758 ;
        RECT 52.342 65.739 57.414 65.804 ;
        RECT 52.296 65.785 57.368 65.85 ;
        RECT 52.25 65.831 57.322 65.896 ;
        RECT 52.204 65.877 57.276 65.942 ;
        RECT 52.158 65.923 57.23 65.988 ;
        RECT 52.112 65.969 57.184 66.034 ;
        RECT 52.066 66.015 57.138 66.08 ;
        RECT 52.02 66.061 57.092 66.126 ;
        RECT 51.974 66.107 57.046 66.172 ;
        RECT 51.928 66.153 57 66.218 ;
        RECT 51.882 66.199 56.954 66.264 ;
        RECT 51.836 66.245 56.908 66.31 ;
        RECT 51.79 66.291 56.862 66.356 ;
        RECT 51.744 66.337 56.816 66.402 ;
        RECT 51.698 66.383 56.77 66.448 ;
        RECT 51.652 66.429 56.724 66.494 ;
        RECT 51.606 66.475 56.678 66.54 ;
        RECT 51.56 66.521 56.632 66.586 ;
        RECT 51.514 66.567 56.586 66.632 ;
        RECT 51.468 66.613 56.54 66.678 ;
        RECT 51.422 66.659 56.494 66.724 ;
        RECT 51.376 66.705 56.448 66.77 ;
        RECT 51.33 66.751 56.402 66.816 ;
        RECT 51.284 66.797 56.356 66.862 ;
        RECT 51.238 66.843 56.31 66.908 ;
        RECT 51.192 66.889 56.264 66.954 ;
        RECT 51.146 66.935 56.218 67 ;
        RECT 51.1 66.981 56.172 67.046 ;
        RECT 51.054 67.027 56.126 67.092 ;
        RECT 51.008 67.073 56.08 67.138 ;
        RECT 50.962 67.119 56.034 67.184 ;
        RECT 50.916 67.165 55.988 67.23 ;
        RECT 50.87 67.211 55.942 67.276 ;
        RECT 50.824 67.257 55.896 67.322 ;
        RECT 50.778 67.303 55.85 67.368 ;
        RECT 50.732 67.349 55.804 67.414 ;
        RECT 50.686 67.395 55.758 67.46 ;
        RECT 50.64 67.441 55.712 67.506 ;
        RECT 50.594 67.487 55.666 67.552 ;
        RECT 50.548 67.533 55.62 67.598 ;
        RECT 50.502 67.579 55.574 67.644 ;
        RECT 50.456 67.625 55.528 67.69 ;
        RECT 50.41 67.671 55.482 67.736 ;
        RECT 50.364 67.717 55.436 67.782 ;
        RECT 50.318 67.763 55.39 67.828 ;
        RECT 50.272 67.809 55.344 67.874 ;
        RECT 50.226 67.855 55.298 67.92 ;
        RECT 50.18 67.901 55.252 67.966 ;
        RECT 50.134 67.947 55.206 68.012 ;
        RECT 50.088 67.993 55.16 68.058 ;
        RECT 50.042 68.039 55.114 68.104 ;
        RECT 49.996 68.085 55.068 68.15 ;
        RECT 49.95 68.131 55.022 68.196 ;
        RECT 49.95 68.131 54.976 68.242 ;
        RECT 49.95 68.131 54.93 68.288 ;
        RECT 49.95 68.131 54.884 68.334 ;
        RECT 49.95 68.131 54.838 68.38 ;
        RECT 49.95 68.131 54.792 68.426 ;
        RECT 49.95 68.131 54.746 68.472 ;
        RECT 49.95 68.131 54.7 68.518 ;
        RECT 49.95 68.131 54.654 68.564 ;
        RECT 49.95 68.131 54.608 68.61 ;
        RECT 49.95 68.131 54.562 68.656 ;
        RECT 49.95 68.131 54.516 68.702 ;
        RECT 49.95 68.131 54.47 68.748 ;
        RECT 49.95 68.131 54.424 68.794 ;
        RECT 49.95 68.131 54.378 68.84 ;
        RECT 49.95 68.131 54.332 68.886 ;
        RECT 49.95 68.131 54.286 68.932 ;
        RECT 49.95 68.131 54.24 68.978 ;
        RECT 49.95 68.131 54.194 69.024 ;
        RECT 49.95 68.131 54.148 69.07 ;
        RECT 49.95 68.131 54.102 69.116 ;
        RECT 49.95 68.131 54.056 69.162 ;
        RECT 49.95 68.131 54.01 69.208 ;
        RECT 49.95 68.131 53.964 69.254 ;
        RECT 49.95 68.131 53.918 69.3 ;
        RECT 49.95 68.131 53.872 69.346 ;
        RECT 49.95 68.131 53.826 69.392 ;
        RECT 49.95 68.131 53.78 69.438 ;
        RECT 49.95 68.131 53.734 69.484 ;
        RECT 49.95 68.131 53.688 69.53 ;
        RECT 49.95 68.131 53.642 69.576 ;
        RECT 49.95 68.131 53.596 69.622 ;
        RECT 49.95 68.131 53.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 54.814 43.323 59.874 43.4 ;
        RECT 59.736 38.401 80 39.45 ;
        RECT 59.828 38.309 59.874 43.4 ;
        RECT 54.768 43.369 59.828 43.446 ;
        RECT 59.782 38.355 80 39.45 ;
        RECT 54.722 43.415 59.782 43.492 ;
        RECT 54.676 43.461 59.736 43.538 ;
        RECT 54.63 43.507 59.69 43.584 ;
        RECT 54.584 43.553 59.644 43.63 ;
        RECT 54.538 43.599 59.598 43.676 ;
        RECT 54.492 43.645 59.552 43.722 ;
        RECT 54.446 43.691 59.506 43.768 ;
        RECT 54.4 43.737 59.46 43.814 ;
        RECT 54.354 43.783 59.414 43.86 ;
        RECT 54.308 43.829 59.368 43.906 ;
        RECT 54.262 43.875 59.322 43.952 ;
        RECT 54.216 43.921 59.276 43.998 ;
        RECT 54.17 43.967 59.23 44.044 ;
        RECT 54.124 44.013 59.184 44.09 ;
        RECT 54.078 44.059 59.138 44.136 ;
        RECT 54.032 44.105 59.092 44.182 ;
        RECT 53.986 44.151 59.046 44.228 ;
        RECT 53.94 44.197 59 44.274 ;
        RECT 53.894 44.243 58.954 44.32 ;
        RECT 53.848 44.289 58.908 44.366 ;
        RECT 53.802 44.335 58.862 44.412 ;
        RECT 53.756 44.381 58.816 44.458 ;
        RECT 53.71 44.427 58.77 44.504 ;
        RECT 53.664 44.473 58.724 44.55 ;
        RECT 53.618 44.519 58.678 44.596 ;
        RECT 53.572 44.565 58.632 44.642 ;
        RECT 53.526 44.611 58.586 44.688 ;
        RECT 53.48 44.657 58.54 44.734 ;
        RECT 53.434 44.703 58.494 44.78 ;
        RECT 53.388 44.749 58.448 44.826 ;
        RECT 53.342 44.795 58.402 44.872 ;
        RECT 53.296 44.841 58.356 44.918 ;
        RECT 53.25 44.887 58.31 44.964 ;
        RECT 53.204 44.933 58.264 45.01 ;
        RECT 53.158 44.979 58.218 45.056 ;
        RECT 53.112 45.025 58.172 45.102 ;
        RECT 53.066 45.071 58.126 45.148 ;
        RECT 53.02 45.117 58.08 45.194 ;
        RECT 52.974 45.163 58.034 45.24 ;
        RECT 52.928 45.209 57.988 45.286 ;
        RECT 52.882 45.255 57.942 45.332 ;
        RECT 52.836 45.301 57.896 45.378 ;
        RECT 52.79 45.347 57.85 45.424 ;
        RECT 52.744 45.393 57.804 45.47 ;
        RECT 52.698 45.439 57.758 45.516 ;
        RECT 52.652 45.485 57.712 45.562 ;
        RECT 52.606 45.531 57.666 45.608 ;
        RECT 52.56 45.577 57.62 45.654 ;
        RECT 52.514 45.623 57.574 45.7 ;
        RECT 52.468 45.669 57.528 45.746 ;
        RECT 52.422 45.715 57.482 45.792 ;
        RECT 52.376 45.761 57.436 45.838 ;
        RECT 52.33 45.807 57.39 45.884 ;
        RECT 52.284 45.853 57.344 45.93 ;
        RECT 52.238 45.899 57.298 45.976 ;
        RECT 52.192 45.945 57.252 46.022 ;
        RECT 52.146 45.991 57.206 46.068 ;
        RECT 52.1 46.037 57.16 46.114 ;
        RECT 52.054 46.083 57.114 46.16 ;
        RECT 52.008 46.129 57.068 46.206 ;
        RECT 51.962 46.175 57.022 46.252 ;
        RECT 51.916 46.221 56.976 46.298 ;
        RECT 51.87 46.267 56.93 46.344 ;
        RECT 51.824 46.313 56.884 46.39 ;
        RECT 51.778 46.359 56.838 46.436 ;
        RECT 51.732 46.405 56.792 46.482 ;
        RECT 51.686 46.451 56.746 46.528 ;
        RECT 51.64 46.497 56.7 46.574 ;
        RECT 51.594 46.543 56.654 46.62 ;
        RECT 51.548 46.589 56.608 46.666 ;
        RECT 51.502 46.635 56.562 46.712 ;
        RECT 51.456 46.681 56.516 46.758 ;
        RECT 51.41 46.727 56.47 46.804 ;
        RECT 51.364 46.773 56.424 46.85 ;
        RECT 51.318 46.819 56.378 46.896 ;
        RECT 51.272 46.865 56.332 46.942 ;
        RECT 51.226 46.911 56.286 46.988 ;
        RECT 51.18 46.957 56.24 47.034 ;
        RECT 51.134 47.003 56.194 47.08 ;
        RECT 51.088 47.049 56.148 47.126 ;
        RECT 51.042 47.095 56.102 47.172 ;
        RECT 50.996 47.141 56.056 47.218 ;
        RECT 50.95 47.187 56.01 47.264 ;
        RECT 50.904 47.233 55.964 47.31 ;
        RECT 50.858 47.279 55.918 47.356 ;
        RECT 50.812 47.325 55.872 47.402 ;
        RECT 50.766 47.371 55.826 47.448 ;
        RECT 50.72 47.417 55.78 47.494 ;
        RECT 50.674 47.463 55.734 47.54 ;
        RECT 50.628 47.509 55.688 47.586 ;
        RECT 50.582 47.555 55.642 47.632 ;
        RECT 50.536 47.601 55.596 47.678 ;
        RECT 50.49 47.647 55.55 47.724 ;
        RECT 50.444 47.693 55.504 47.77 ;
        RECT 50.398 47.739 55.458 47.816 ;
        RECT 50.352 47.785 55.412 47.862 ;
        RECT 50.306 47.831 55.366 47.908 ;
        RECT 50.26 47.877 55.32 47.954 ;
        RECT 50.214 47.923 55.274 48 ;
        RECT 50.168 47.969 55.228 48.046 ;
        RECT 50.122 48.015 55.182 48.092 ;
        RECT 50.076 48.061 55.136 48.138 ;
        RECT 50.03 48.107 55.09 48.184 ;
        RECT 49.984 48.153 55.044 48.23 ;
        RECT 49.938 48.199 54.998 48.276 ;
        RECT 49.892 48.245 54.952 48.322 ;
        RECT 49.846 48.291 54.906 48.368 ;
        RECT 49.8 48.337 54.86 48.414 ;
        RECT 49.754 48.383 54.814 48.46 ;
        RECT 49.708 48.429 54.768 48.506 ;
        RECT 49.662 48.475 54.722 48.552 ;
        RECT 49.616 48.521 54.676 48.598 ;
        RECT 49.57 48.567 54.63 48.644 ;
        RECT 49.524 48.613 54.584 48.69 ;
        RECT 49.478 48.659 54.538 48.736 ;
        RECT 49.432 48.705 54.492 48.782 ;
        RECT 49.386 48.751 54.446 48.828 ;
        RECT 49.34 48.797 54.4 48.874 ;
        RECT 49.294 48.843 54.354 48.92 ;
        RECT 49.248 48.889 54.308 48.966 ;
        RECT 49.202 48.935 54.262 49.012 ;
        RECT 49.156 48.981 54.216 49.058 ;
        RECT 49.11 49.027 54.17 49.104 ;
        RECT 49.064 49.073 54.124 49.15 ;
        RECT 49.018 49.119 54.078 49.196 ;
        RECT 48.972 49.165 54.032 49.242 ;
        RECT 48.926 49.211 53.986 49.288 ;
        RECT 48.88 49.257 53.94 49.334 ;
        RECT 48.834 49.303 53.894 49.38 ;
        RECT 48.788 49.349 53.848 49.426 ;
        RECT 48.742 49.395 53.802 49.472 ;
        RECT 48.696 49.441 53.756 49.518 ;
        RECT 48.65 49.487 53.71 49.564 ;
        RECT 48.604 49.533 53.664 49.61 ;
        RECT 48.558 49.579 53.618 49.656 ;
        RECT 48.512 49.625 53.572 49.702 ;
        RECT 48.466 49.671 53.526 49.748 ;
        RECT 48.42 49.717 53.48 49.794 ;
        RECT 48.374 49.763 53.434 49.84 ;
        RECT 48.328 49.809 53.388 49.886 ;
        RECT 48.282 49.855 53.342 49.932 ;
        RECT 48.236 49.901 53.296 49.978 ;
        RECT 48.19 49.947 53.25 50.024 ;
        RECT 48.144 49.993 53.204 50.07 ;
        RECT 48.098 50.039 53.158 50.116 ;
        RECT 48.052 50.085 53.112 50.162 ;
        RECT 48.006 50.131 53.066 50.208 ;
        RECT 47.96 50.177 53.02 50.254 ;
        RECT 47.914 50.223 52.974 50.3 ;
        RECT 47.868 50.269 52.928 50.346 ;
        RECT 47.822 50.315 52.882 50.392 ;
        RECT 47.776 50.361 52.836 50.438 ;
        RECT 47.73 50.407 52.79 50.484 ;
        RECT 47.684 50.453 52.744 50.53 ;
        RECT 47.638 50.499 52.698 50.576 ;
        RECT 47.592 50.545 52.652 50.622 ;
        RECT 47.546 50.591 52.606 50.668 ;
        RECT 47.5 50.637 52.56 50.714 ;
        RECT 47.454 50.683 52.514 50.76 ;
        RECT 47.408 50.729 52.468 50.806 ;
        RECT 47.362 50.775 52.422 50.852 ;
        RECT 47.316 50.821 52.376 50.898 ;
        RECT 47.27 50.867 52.33 50.944 ;
        RECT 47.224 50.913 52.284 50.99 ;
        RECT 47.178 50.959 52.238 51.036 ;
        RECT 47.132 51.005 52.192 51.082 ;
        RECT 47.086 51.051 52.146 51.128 ;
        RECT 47.04 51.097 52.1 51.174 ;
        RECT 46.994 51.143 52.054 51.22 ;
        RECT 46.948 51.189 52.008 51.266 ;
        RECT 46.902 51.235 51.962 51.312 ;
        RECT 46.856 51.281 51.916 51.358 ;
        RECT 46.81 51.327 51.87 51.404 ;
        RECT 46.764 51.373 51.824 51.45 ;
        RECT 46.718 51.419 51.778 51.496 ;
        RECT 46.672 51.465 51.732 51.542 ;
        RECT 46.626 51.511 51.686 51.588 ;
        RECT 46.58 51.557 51.64 51.634 ;
        RECT 46.534 51.603 51.594 51.68 ;
        RECT 46.488 51.649 51.548 51.726 ;
        RECT 46.442 51.695 51.502 51.772 ;
        RECT 46.396 51.741 51.456 51.818 ;
        RECT 46.35 51.787 51.41 51.864 ;
        RECT 46.304 51.833 51.364 51.91 ;
        RECT 46.258 51.879 51.318 51.956 ;
        RECT 46.212 51.925 51.272 52.002 ;
        RECT 46.166 51.971 51.226 52.048 ;
        RECT 46.12 52.017 51.18 52.094 ;
        RECT 46.074 52.063 51.134 52.14 ;
        RECT 46.028 52.109 51.088 52.186 ;
        RECT 45.982 52.155 51.042 52.232 ;
        RECT 45.936 52.201 50.996 52.278 ;
        RECT 45.89 52.247 50.95 52.324 ;
        RECT 45.844 52.293 50.904 52.37 ;
        RECT 45.798 52.339 50.858 52.416 ;
        RECT 45.752 52.385 50.812 52.462 ;
        RECT 45.706 52.431 50.766 52.508 ;
        RECT 45.66 52.477 50.72 52.554 ;
        RECT 45.614 52.523 50.674 52.6 ;
        RECT 45.568 52.569 50.628 52.646 ;
        RECT 45.522 52.615 50.582 52.692 ;
        RECT 45.476 52.661 50.536 52.738 ;
        RECT 45.43 52.707 50.49 52.784 ;
        RECT 45.384 52.753 50.444 52.83 ;
        RECT 45.338 52.799 50.398 52.876 ;
        RECT 45.292 52.845 50.352 52.922 ;
        RECT 45.246 52.891 50.306 52.968 ;
        RECT 45.2 52.937 50.26 53.014 ;
        RECT 45.154 52.983 50.214 53.06 ;
        RECT 45.108 53.029 50.168 53.106 ;
        RECT 45.062 53.075 50.122 53.152 ;
        RECT 45.016 53.121 50.076 53.198 ;
        RECT 44.97 53.167 50.03 53.244 ;
        RECT 44.924 53.213 49.984 53.29 ;
        RECT 44.878 53.259 49.938 53.336 ;
        RECT 44.832 53.305 49.892 53.382 ;
        RECT 44.786 53.351 49.846 53.428 ;
        RECT 44.74 53.397 49.8 53.474 ;
        RECT 44.694 53.443 49.754 53.52 ;
        RECT 44.648 53.489 49.708 53.566 ;
        RECT 44.602 53.535 49.662 53.612 ;
        RECT 44.556 53.581 49.616 53.658 ;
        RECT 44.51 53.627 49.57 53.704 ;
        RECT 44.464 53.673 49.524 53.75 ;
        RECT 44.418 53.719 49.478 53.796 ;
        RECT 44.372 53.765 49.432 53.842 ;
        RECT 44.326 53.811 49.386 53.888 ;
        RECT 44.28 53.857 49.34 53.934 ;
        RECT 44.234 53.903 49.294 53.98 ;
        RECT 44.188 53.949 49.248 54.026 ;
        RECT 44.142 53.995 49.202 54.072 ;
        RECT 44.096 54.041 49.156 54.118 ;
        RECT 44.05 54.087 49.11 54.164 ;
        RECT 44.004 54.133 49.064 54.21 ;
        RECT 43.958 54.179 49.018 54.256 ;
        RECT 43.912 54.225 48.972 54.302 ;
        RECT 43.866 54.271 48.926 54.348 ;
        RECT 43.82 54.317 48.88 54.394 ;
        RECT 43.774 54.363 48.834 54.44 ;
        RECT 43.728 54.409 48.788 54.486 ;
        RECT 43.682 54.455 48.742 54.532 ;
        RECT 43.636 54.501 48.696 54.578 ;
        RECT 43.59 54.547 48.65 54.624 ;
        RECT 43.544 54.593 48.604 54.67 ;
        RECT 43.498 54.639 48.558 54.716 ;
        RECT 43.452 54.685 48.512 54.762 ;
        RECT 43.406 54.731 48.466 54.808 ;
        RECT 43.36 54.777 48.42 54.854 ;
        RECT 43.314 54.823 48.374 54.9 ;
        RECT 43.268 54.869 48.328 54.946 ;
        RECT 43.222 54.915 48.282 54.992 ;
        RECT 43.176 54.961 48.236 55.038 ;
        RECT 43.13 55.007 48.19 55.084 ;
        RECT 43.084 55.053 48.144 55.13 ;
        RECT 43.038 55.099 48.098 55.176 ;
        RECT 42.992 55.145 48.052 55.222 ;
        RECT 42.946 55.191 48.006 55.268 ;
        RECT 42.9 55.237 47.96 55.314 ;
        RECT 42.854 55.283 47.914 55.36 ;
        RECT 42.808 55.329 47.868 55.406 ;
        RECT 42.762 55.375 47.822 55.452 ;
        RECT 42.716 55.421 47.776 55.498 ;
        RECT 42.67 55.467 47.73 55.544 ;
        RECT 42.624 55.513 47.684 55.59 ;
        RECT 42.578 55.559 47.638 55.636 ;
        RECT 42.532 55.605 47.592 55.682 ;
        RECT 42.486 55.651 47.546 55.728 ;
        RECT 42.44 55.697 47.5 55.774 ;
        RECT 42.394 55.743 47.454 55.82 ;
        RECT 42.348 55.789 47.408 55.866 ;
        RECT 42.302 55.835 47.362 55.912 ;
        RECT 42.256 55.881 47.316 55.958 ;
        RECT 42.21 55.927 47.27 56.004 ;
        RECT 42.164 55.973 47.224 56.05 ;
        RECT 42.118 56.019 47.178 56.096 ;
        RECT 42.072 56.065 47.132 56.142 ;
        RECT 42.026 56.111 47.086 56.188 ;
        RECT 41.98 56.157 47.04 56.234 ;
        RECT 41.934 56.203 46.994 56.28 ;
        RECT 41.888 56.249 46.948 56.326 ;
        RECT 41.842 56.295 46.902 56.372 ;
        RECT 41.796 56.341 46.856 56.418 ;
        RECT 41.75 56.387 46.81 56.464 ;
        RECT 41.704 56.433 46.764 56.51 ;
        RECT 41.658 56.479 46.718 56.556 ;
        RECT 41.612 56.525 46.672 56.602 ;
        RECT 41.566 56.571 46.626 56.648 ;
        RECT 41.52 56.617 46.58 56.694 ;
        RECT 41.474 56.663 46.534 56.74 ;
        RECT 41.428 56.709 46.488 56.786 ;
        RECT 41.382 56.755 46.442 56.832 ;
        RECT 41.336 56.801 46.396 56.878 ;
        RECT 41.29 56.847 46.35 56.924 ;
        RECT 41.244 56.893 46.304 56.97 ;
        RECT 41.198 56.939 46.258 57.016 ;
        RECT 41.152 56.985 46.212 57.062 ;
        RECT 41.106 57.031 46.166 57.108 ;
        RECT 41.06 57.077 46.12 57.154 ;
        RECT 41.014 57.123 46.074 57.2 ;
        RECT 40.968 57.169 46.028 57.246 ;
        RECT 40.922 57.215 45.982 57.292 ;
        RECT 40.876 57.261 45.936 57.338 ;
        RECT 40.83 57.307 45.89 57.384 ;
        RECT 40.784 57.353 45.844 57.43 ;
        RECT 40.738 57.399 45.798 57.476 ;
        RECT 40.692 57.445 45.752 57.522 ;
        RECT 40.646 57.491 45.706 57.568 ;
        RECT 40.6 57.537 45.66 57.614 ;
        RECT 40.554 57.583 45.614 57.66 ;
        RECT 40.508 57.629 45.568 57.706 ;
        RECT 40.462 57.675 45.522 57.752 ;
        RECT 40.416 57.721 45.476 57.798 ;
        RECT 40.37 57.767 45.43 57.844 ;
        RECT 40.324 57.813 45.384 57.89 ;
        RECT 40.278 57.859 45.338 57.936 ;
        RECT 40.232 57.905 45.292 57.982 ;
        RECT 40.186 57.951 45.246 58.028 ;
        RECT 40.14 57.997 45.2 58.074 ;
        RECT 40.094 58.043 45.154 58.12 ;
        RECT 40.048 58.089 45.108 58.166 ;
        RECT 40.002 58.135 45.062 58.212 ;
        RECT 39.956 58.181 45.016 58.258 ;
        RECT 39.91 58.227 44.97 58.304 ;
        RECT 39.864 58.273 44.924 58.35 ;
        RECT 39.818 58.319 44.878 58.396 ;
        RECT 39.772 58.365 44.832 58.442 ;
        RECT 39.726 58.411 44.786 58.488 ;
        RECT 39.68 58.457 44.74 58.534 ;
        RECT 39.634 58.503 44.694 58.58 ;
        RECT 39.588 58.549 44.648 58.626 ;
        RECT 39.542 58.595 44.602 58.672 ;
        RECT 39.45 58.687 44.556 58.718 ;
        RECT 39.496 58.641 44.556 58.718 ;
        RECT 39.438 58.716 44.51 58.764 ;
        RECT 39.392 58.745 44.464 58.81 ;
        RECT 39.346 58.791 44.418 58.856 ;
        RECT 39.3 58.837 44.372 58.902 ;
        RECT 39.254 58.883 44.326 58.948 ;
        RECT 39.208 58.929 44.28 58.994 ;
        RECT 39.162 58.975 44.234 59.04 ;
        RECT 39.116 59.021 44.188 59.086 ;
        RECT 39.07 59.067 44.142 59.132 ;
        RECT 39.024 59.113 44.096 59.178 ;
        RECT 38.978 59.159 44.05 59.224 ;
        RECT 38.932 59.205 44.004 59.27 ;
        RECT 38.886 59.251 43.958 59.316 ;
        RECT 38.84 59.297 43.912 59.362 ;
        RECT 38.794 59.343 43.866 59.408 ;
        RECT 38.748 59.389 43.82 59.454 ;
        RECT 38.702 59.435 43.774 59.5 ;
        RECT 38.656 59.481 43.728 59.546 ;
        RECT 38.61 59.527 43.682 59.592 ;
        RECT 38.564 59.573 43.636 59.638 ;
        RECT 38.518 59.619 43.59 59.684 ;
        RECT 38.472 59.665 43.544 59.73 ;
        RECT 38.426 59.711 43.498 59.776 ;
        RECT 38.38 59.757 43.452 59.822 ;
        RECT 38.334 59.803 43.406 59.868 ;
        RECT 38.288 59.849 43.36 59.914 ;
        RECT 38.242 59.895 43.314 59.96 ;
        RECT 38.196 59.941 43.268 60.006 ;
        RECT 38.15 59.987 43.222 60.052 ;
        RECT 38.104 60.033 43.176 60.098 ;
        RECT 38.058 60.079 43.13 60.144 ;
        RECT 38.012 60.125 43.084 60.19 ;
        RECT 37.966 60.171 43.038 60.236 ;
        RECT 37.92 60.217 42.992 60.282 ;
        RECT 37.874 60.263 42.946 60.328 ;
        RECT 37.828 60.309 42.9 60.374 ;
        RECT 37.782 60.355 42.854 60.42 ;
        RECT 37.736 60.401 42.808 60.466 ;
        RECT 37.69 60.447 42.762 60.512 ;
        RECT 37.644 60.493 42.716 60.558 ;
        RECT 37.598 60.539 42.67 60.604 ;
        RECT 37.552 60.585 42.624 60.65 ;
        RECT 37.506 60.631 42.578 60.696 ;
        RECT 37.46 60.677 42.532 60.742 ;
        RECT 37.414 60.723 42.486 60.788 ;
        RECT 37.368 60.769 42.44 60.834 ;
        RECT 37.322 60.815 42.394 60.88 ;
        RECT 37.276 60.861 42.348 60.926 ;
        RECT 37.23 60.907 42.302 60.972 ;
        RECT 37.184 60.953 42.256 61.018 ;
        RECT 37.138 60.999 42.21 61.064 ;
        RECT 37.092 61.045 42.164 61.11 ;
        RECT 37.046 61.091 42.118 61.156 ;
        RECT 37 61.137 42.072 61.202 ;
        RECT 36.954 61.183 42.026 61.248 ;
        RECT 36.908 61.229 41.98 61.294 ;
        RECT 36.862 61.275 41.934 61.34 ;
        RECT 36.816 61.321 41.888 61.386 ;
        RECT 36.77 61.367 41.842 61.432 ;
        RECT 36.724 61.413 41.796 61.478 ;
        RECT 36.678 61.459 41.75 61.524 ;
        RECT 36.632 61.505 41.704 61.57 ;
        RECT 36.586 61.551 41.658 61.616 ;
        RECT 36.54 61.597 41.612 61.662 ;
        RECT 36.494 61.643 41.566 61.708 ;
        RECT 36.448 61.689 41.52 61.754 ;
        RECT 36.402 61.735 41.474 61.8 ;
        RECT 36.356 61.781 41.428 61.846 ;
        RECT 36.31 61.827 41.382 61.892 ;
        RECT 36.264 61.873 41.336 61.938 ;
        RECT 36.218 61.919 41.29 61.984 ;
        RECT 36.172 61.965 41.244 62.03 ;
        RECT 36.126 62.011 41.198 62.076 ;
        RECT 36.08 62.057 41.152 62.122 ;
        RECT 36.034 62.103 41.106 62.168 ;
        RECT 35.988 62.149 41.06 62.214 ;
        RECT 35.942 62.195 41.014 62.26 ;
        RECT 35.896 62.241 40.968 62.306 ;
        RECT 35.85 62.287 40.922 62.352 ;
        RECT 35.85 62.287 40.876 62.398 ;
        RECT 35.85 62.287 40.83 62.444 ;
        RECT 35.85 62.287 40.784 62.49 ;
        RECT 35.85 62.287 40.738 62.536 ;
        RECT 35.85 62.287 40.692 62.582 ;
        RECT 35.85 62.287 40.646 62.628 ;
        RECT 35.85 62.287 40.6 62.674 ;
        RECT 35.85 62.287 40.554 62.72 ;
        RECT 35.85 62.287 40.508 62.766 ;
        RECT 35.85 62.287 40.462 62.812 ;
        RECT 35.85 62.287 40.416 62.858 ;
        RECT 35.85 62.287 40.37 62.904 ;
        RECT 35.85 62.287 40.324 62.95 ;
        RECT 35.85 62.287 40.278 62.996 ;
        RECT 35.85 62.287 40.232 63.042 ;
        RECT 35.85 62.287 40.186 63.088 ;
        RECT 35.85 62.287 40.14 63.134 ;
        RECT 35.85 62.287 40.094 63.18 ;
        RECT 35.85 62.287 40.048 63.226 ;
        RECT 35.85 62.287 40.002 63.272 ;
        RECT 35.85 62.287 39.956 63.318 ;
        RECT 35.85 62.287 39.91 63.364 ;
        RECT 35.85 62.287 39.864 63.41 ;
        RECT 35.85 62.287 39.818 63.456 ;
        RECT 35.85 62.287 39.772 63.502 ;
        RECT 35.85 62.287 39.726 63.548 ;
        RECT 35.85 62.287 39.68 63.594 ;
        RECT 35.85 62.287 39.634 63.64 ;
        RECT 35.85 62.287 39.588 63.686 ;
        RECT 35.85 62.287 39.542 63.732 ;
        RECT 35.85 62.287 39.496 63.778 ;
        RECT 35.85 62.287 39.45 80 ;
        RECT 62.31 35.85 80 39.45 ;
        RECT 58.678 39.459 63.782 39.492 ;
        RECT 57.252 40.885 62.31 40.963 ;
        RECT 57.298 40.839 62.356 40.918 ;
        RECT 62.266 35.872 62.31 40.963 ;
        RECT 57.206 40.931 62.266 41.008 ;
        RECT 57.344 40.793 62.402 40.872 ;
        RECT 62.22 35.917 62.266 41.008 ;
        RECT 57.16 40.977 62.22 41.054 ;
        RECT 57.39 40.747 62.448 40.826 ;
        RECT 62.174 35.963 62.22 41.054 ;
        RECT 57.114 41.023 62.174 41.1 ;
        RECT 57.436 40.701 62.494 40.78 ;
        RECT 62.128 36.009 62.174 41.1 ;
        RECT 57.068 41.069 62.128 41.146 ;
        RECT 57.482 40.655 62.54 40.734 ;
        RECT 62.082 36.055 62.128 41.146 ;
        RECT 57.022 41.115 62.082 41.192 ;
        RECT 57.528 40.609 62.586 40.688 ;
        RECT 62.036 36.101 62.082 41.192 ;
        RECT 56.976 41.161 62.036 41.238 ;
        RECT 57.574 40.563 62.632 40.642 ;
        RECT 61.99 36.147 62.036 41.238 ;
        RECT 56.93 41.207 61.99 41.284 ;
        RECT 57.62 40.517 62.678 40.596 ;
        RECT 61.944 36.193 61.99 41.284 ;
        RECT 56.884 41.253 61.944 41.33 ;
        RECT 57.666 40.471 62.724 40.55 ;
        RECT 61.898 36.239 61.944 41.33 ;
        RECT 56.838 41.299 61.898 41.376 ;
        RECT 57.712 40.425 62.77 40.504 ;
        RECT 61.852 36.285 61.898 41.376 ;
        RECT 56.792 41.345 61.852 41.422 ;
        RECT 57.758 40.379 62.816 40.458 ;
        RECT 61.806 36.331 61.852 41.422 ;
        RECT 56.746 41.391 61.806 41.468 ;
        RECT 57.804 40.333 62.862 40.412 ;
        RECT 61.76 36.377 61.806 41.468 ;
        RECT 56.7 41.437 61.76 41.514 ;
        RECT 57.85 40.287 62.908 40.366 ;
        RECT 61.714 36.423 61.76 41.514 ;
        RECT 56.654 41.483 61.714 41.56 ;
        RECT 57.896 40.241 62.954 40.32 ;
        RECT 61.668 36.469 61.714 41.56 ;
        RECT 56.608 41.529 61.668 41.606 ;
        RECT 57.942 40.195 63 40.274 ;
        RECT 61.622 36.515 61.668 41.606 ;
        RECT 56.562 41.575 61.622 41.652 ;
        RECT 57.988 40.149 63.046 40.228 ;
        RECT 61.576 36.561 61.622 41.652 ;
        RECT 56.516 41.621 61.576 41.698 ;
        RECT 58.034 40.103 63.092 40.182 ;
        RECT 61.53 36.607 61.576 41.698 ;
        RECT 56.47 41.667 61.53 41.744 ;
        RECT 58.08 40.057 63.138 40.136 ;
        RECT 61.484 36.653 61.53 41.744 ;
        RECT 56.424 41.713 61.484 41.79 ;
        RECT 58.126 40.011 63.184 40.09 ;
        RECT 61.438 36.699 61.484 41.79 ;
        RECT 56.378 41.759 61.438 41.836 ;
        RECT 58.172 39.965 63.23 40.044 ;
        RECT 61.392 36.745 61.438 41.836 ;
        RECT 56.332 41.805 61.392 41.882 ;
        RECT 58.218 39.919 63.276 39.998 ;
        RECT 61.346 36.791 61.392 41.882 ;
        RECT 56.286 41.851 61.346 41.928 ;
        RECT 58.264 39.873 63.322 39.952 ;
        RECT 61.3 36.837 61.346 41.928 ;
        RECT 56.24 41.897 61.3 41.974 ;
        RECT 58.31 39.827 63.368 39.906 ;
        RECT 61.254 36.883 61.3 41.974 ;
        RECT 56.194 41.943 61.254 42.02 ;
        RECT 58.356 39.781 63.414 39.86 ;
        RECT 61.208 36.929 61.254 42.02 ;
        RECT 56.148 41.989 61.208 42.066 ;
        RECT 58.402 39.735 63.46 39.814 ;
        RECT 61.162 36.975 61.208 42.066 ;
        RECT 56.102 42.035 61.162 42.112 ;
        RECT 58.448 39.689 63.506 39.768 ;
        RECT 61.116 37.021 61.162 42.112 ;
        RECT 56.056 42.081 61.116 42.158 ;
        RECT 58.494 39.643 63.552 39.722 ;
        RECT 61.07 37.067 61.116 42.158 ;
        RECT 56.01 42.127 61.07 42.204 ;
        RECT 58.54 39.597 63.598 39.676 ;
        RECT 61.024 37.113 61.07 42.204 ;
        RECT 55.964 42.173 61.024 42.25 ;
        RECT 58.586 39.551 63.644 39.63 ;
        RECT 60.978 37.159 61.024 42.25 ;
        RECT 55.918 42.219 60.978 42.296 ;
        RECT 58.632 39.505 63.69 39.584 ;
        RECT 60.932 37.205 60.978 42.296 ;
        RECT 55.872 42.265 60.932 42.342 ;
        RECT 58.678 39.459 63.736 39.538 ;
        RECT 60.886 37.251 60.932 42.342 ;
        RECT 55.826 42.311 60.886 42.388 ;
        RECT 58.724 39.413 63.801 39.46 ;
        RECT 60.84 37.297 60.886 42.388 ;
        RECT 55.78 42.357 60.84 42.434 ;
        RECT 58.77 39.367 80 39.45 ;
        RECT 60.794 37.343 60.84 42.434 ;
        RECT 55.734 42.403 60.794 42.48 ;
        RECT 58.816 39.321 80 39.45 ;
        RECT 60.748 37.389 60.794 42.48 ;
        RECT 55.688 42.449 60.748 42.526 ;
        RECT 58.862 39.275 80 39.45 ;
        RECT 60.702 37.435 60.748 42.526 ;
        RECT 55.642 42.495 60.702 42.572 ;
        RECT 58.908 39.229 80 39.45 ;
        RECT 60.656 37.481 60.702 42.572 ;
        RECT 55.596 42.541 60.656 42.618 ;
        RECT 58.954 39.183 80 39.45 ;
        RECT 60.61 37.527 60.656 42.618 ;
        RECT 55.55 42.587 60.61 42.664 ;
        RECT 59 39.137 80 39.45 ;
        RECT 60.564 37.573 60.61 42.664 ;
        RECT 55.504 42.633 60.564 42.71 ;
        RECT 59.046 39.091 80 39.45 ;
        RECT 60.518 37.619 60.564 42.71 ;
        RECT 55.458 42.679 60.518 42.756 ;
        RECT 59.092 39.045 80 39.45 ;
        RECT 60.472 37.665 60.518 42.756 ;
        RECT 55.412 42.725 60.472 42.802 ;
        RECT 59.138 38.999 80 39.45 ;
        RECT 60.426 37.711 60.472 42.802 ;
        RECT 55.366 42.771 60.426 42.848 ;
        RECT 59.184 38.953 80 39.45 ;
        RECT 60.38 37.757 60.426 42.848 ;
        RECT 55.32 42.817 60.38 42.894 ;
        RECT 59.23 38.907 80 39.45 ;
        RECT 60.334 37.803 60.38 42.894 ;
        RECT 55.274 42.863 60.334 42.94 ;
        RECT 59.276 38.861 80 39.45 ;
        RECT 60.288 37.849 60.334 42.94 ;
        RECT 55.228 42.909 60.288 42.986 ;
        RECT 59.322 38.815 80 39.45 ;
        RECT 60.242 37.895 60.288 42.986 ;
        RECT 55.182 42.955 60.242 43.032 ;
        RECT 59.368 38.769 80 39.45 ;
        RECT 60.196 37.941 60.242 43.032 ;
        RECT 55.136 43.001 60.196 43.078 ;
        RECT 59.414 38.723 80 39.45 ;
        RECT 60.15 37.987 60.196 43.078 ;
        RECT 55.09 43.047 60.15 43.124 ;
        RECT 59.46 38.677 80 39.45 ;
        RECT 60.104 38.033 60.15 43.124 ;
        RECT 55.044 43.093 60.104 43.17 ;
        RECT 59.506 38.631 80 39.45 ;
        RECT 60.058 38.079 60.104 43.17 ;
        RECT 54.998 43.139 60.058 43.216 ;
        RECT 59.552 38.585 80 39.45 ;
        RECT 60.012 38.125 60.058 43.216 ;
        RECT 54.952 43.185 60.012 43.262 ;
        RECT 59.598 38.539 80 39.45 ;
        RECT 59.966 38.171 60.012 43.262 ;
        RECT 54.906 43.231 59.966 43.308 ;
        RECT 59.644 38.493 80 39.45 ;
        RECT 59.92 38.217 59.966 43.308 ;
        RECT 54.86 43.277 59.92 43.354 ;
        RECT 59.69 38.447 80 39.45 ;
        RECT 59.874 38.263 59.92 43.354 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 77.892 73.45 80 77.05 ;
        RECT 74.278 77.041 79.384 77.06 ;
        RECT 73.45 77.869 78.536 77.921 ;
        RECT 73.45 77.869 78.49 77.967 ;
        RECT 73.45 77.869 78.444 78.013 ;
        RECT 73.45 77.869 78.398 78.059 ;
        RECT 73.45 77.869 78.352 78.105 ;
        RECT 73.45 77.869 78.306 78.151 ;
        RECT 73.45 77.869 78.26 78.197 ;
        RECT 73.45 77.869 78.214 78.243 ;
        RECT 73.45 77.869 78.168 78.289 ;
        RECT 73.45 77.869 78.122 78.335 ;
        RECT 73.45 77.869 78.076 78.381 ;
        RECT 73.45 77.869 78.03 78.427 ;
        RECT 73.45 77.869 77.984 78.473 ;
        RECT 73.45 77.869 77.938 78.519 ;
        RECT 73.496 77.823 78.582 77.875 ;
        RECT 77.878 73.457 77.892 78.549 ;
        RECT 73.542 77.777 78.628 77.829 ;
        RECT 77.832 73.487 77.878 78.579 ;
        RECT 73.588 77.731 78.674 77.783 ;
        RECT 77.786 73.533 77.832 78.625 ;
        RECT 73.634 77.685 78.72 77.737 ;
        RECT 77.74 73.579 77.786 78.671 ;
        RECT 73.68 77.639 78.766 77.691 ;
        RECT 77.694 73.625 77.74 78.717 ;
        RECT 73.726 77.593 78.812 77.645 ;
        RECT 77.648 73.671 77.694 78.763 ;
        RECT 73.772 77.547 78.858 77.599 ;
        RECT 77.602 73.717 77.648 78.809 ;
        RECT 73.818 77.501 78.904 77.553 ;
        RECT 77.556 73.763 77.602 78.855 ;
        RECT 73.864 77.455 78.95 77.507 ;
        RECT 77.51 73.809 77.556 78.901 ;
        RECT 73.91 77.409 78.996 77.461 ;
        RECT 77.464 73.855 77.51 78.947 ;
        RECT 73.956 77.363 79.042 77.415 ;
        RECT 77.418 73.901 77.464 78.993 ;
        RECT 74.002 77.317 79.088 77.369 ;
        RECT 77.372 73.947 77.418 79.039 ;
        RECT 74.048 77.271 79.134 77.323 ;
        RECT 77.326 73.993 77.372 79.085 ;
        RECT 74.094 77.225 79.18 77.277 ;
        RECT 77.28 74.039 77.326 79.131 ;
        RECT 74.14 77.179 79.226 77.231 ;
        RECT 77.234 74.085 77.28 79.177 ;
        RECT 74.186 77.133 79.272 77.185 ;
        RECT 77.188 74.131 77.234 79.223 ;
        RECT 74.232 77.087 79.318 77.139 ;
        RECT 77.142 74.177 77.188 79.269 ;
        RECT 74.278 77.041 79.364 77.093 ;
        RECT 77.096 74.223 77.142 79.315 ;
        RECT 74.324 76.995 80 77.05 ;
        RECT 77.05 74.269 77.096 79.361 ;
        RECT 73.45 77.869 77.05 80 ;
        RECT 74.37 76.949 80 77.05 ;
        RECT 77.038 74.298 77.05 80 ;
        RECT 74.416 76.903 80 77.05 ;
        RECT 76.992 74.327 77.05 80 ;
        RECT 74.462 76.857 80 77.05 ;
        RECT 76.946 74.373 77.05 80 ;
        RECT 74.508 76.811 80 77.05 ;
        RECT 76.9 74.419 77.05 80 ;
        RECT 74.554 76.765 80 77.05 ;
        RECT 76.854 74.465 77.05 80 ;
        RECT 74.6 76.719 80 77.05 ;
        RECT 76.808 74.511 77.05 80 ;
        RECT 74.646 76.673 80 77.05 ;
        RECT 76.762 74.557 77.05 80 ;
        RECT 74.692 76.627 80 77.05 ;
        RECT 76.716 74.603 77.05 80 ;
        RECT 74.738 76.581 80 77.05 ;
        RECT 76.67 74.649 77.05 80 ;
        RECT 74.784 76.535 80 77.05 ;
        RECT 76.624 74.695 77.05 80 ;
        RECT 74.83 76.489 80 77.05 ;
        RECT 76.578 74.741 77.05 80 ;
        RECT 74.876 76.443 80 77.05 ;
        RECT 76.532 74.787 77.05 80 ;
        RECT 74.922 76.397 80 77.05 ;
        RECT 76.486 74.833 77.05 80 ;
        RECT 74.968 76.351 80 77.05 ;
        RECT 76.44 74.879 77.05 80 ;
        RECT 75.014 76.305 80 77.05 ;
        RECT 76.394 74.925 77.05 80 ;
        RECT 75.06 76.259 80 77.05 ;
        RECT 76.348 74.971 77.05 80 ;
        RECT 75.106 76.213 80 77.05 ;
        RECT 76.302 75.017 77.05 80 ;
        RECT 75.152 76.167 80 77.05 ;
        RECT 76.256 75.063 77.05 80 ;
        RECT 75.198 76.121 80 77.05 ;
        RECT 76.21 75.109 77.05 80 ;
        RECT 75.244 76.075 80 77.05 ;
        RECT 76.164 75.155 77.05 80 ;
        RECT 75.29 76.029 80 77.05 ;
        RECT 76.118 75.201 77.05 80 ;
        RECT 75.336 75.983 80 77.05 ;
        RECT 76.072 75.247 77.05 80 ;
        RECT 75.382 75.937 80 77.05 ;
        RECT 76.026 75.293 77.05 80 ;
        RECT 75.428 75.891 80 77.05 ;
        RECT 75.98 75.339 77.05 80 ;
        RECT 75.474 75.845 80 77.05 ;
        RECT 75.934 75.385 77.05 80 ;
        RECT 75.52 75.799 80 77.05 ;
        RECT 75.888 75.431 77.05 80 ;
        RECT 75.566 75.753 80 77.05 ;
        RECT 75.842 75.477 77.05 80 ;
        RECT 75.612 75.707 80 77.05 ;
        RECT 75.796 75.523 77.05 80 ;
        RECT 75.658 75.661 80 77.05 ;
        RECT 75.75 75.569 77.05 80 ;
        RECT 75.704 75.615 80 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 72.05 59.35 80 62.95 ;
        RECT 68.424 62.953 73.522 62.992 ;
        RECT 66.998 64.379 72.05 64.46 ;
        RECT 67.044 64.333 72.096 64.418 ;
        RECT 72.012 59.369 72.05 64.46 ;
        RECT 66.952 64.425 72.012 64.502 ;
        RECT 67.09 64.287 72.142 64.372 ;
        RECT 71.966 59.411 72.012 64.502 ;
        RECT 66.906 64.471 71.966 64.548 ;
        RECT 67.136 64.241 72.188 64.326 ;
        RECT 71.92 59.457 71.966 64.548 ;
        RECT 66.86 64.517 71.92 64.594 ;
        RECT 67.182 64.195 72.234 64.28 ;
        RECT 71.874 59.503 71.92 64.594 ;
        RECT 66.814 64.563 71.874 64.64 ;
        RECT 67.228 64.149 72.28 64.234 ;
        RECT 71.828 59.549 71.874 64.64 ;
        RECT 66.768 64.609 71.828 64.686 ;
        RECT 67.274 64.103 72.326 64.188 ;
        RECT 71.782 59.595 71.828 64.686 ;
        RECT 66.722 64.655 71.782 64.732 ;
        RECT 67.32 64.057 72.372 64.142 ;
        RECT 71.736 59.641 71.782 64.732 ;
        RECT 66.676 64.701 71.736 64.778 ;
        RECT 67.366 64.011 72.418 64.096 ;
        RECT 71.69 59.687 71.736 64.778 ;
        RECT 66.63 64.747 71.69 64.824 ;
        RECT 67.412 63.965 72.464 64.05 ;
        RECT 71.644 59.733 71.69 64.824 ;
        RECT 66.584 64.793 71.644 64.87 ;
        RECT 67.458 63.919 72.51 64.004 ;
        RECT 71.598 59.779 71.644 64.87 ;
        RECT 66.538 64.839 71.598 64.916 ;
        RECT 67.504 63.873 72.556 63.958 ;
        RECT 71.552 59.825 71.598 64.916 ;
        RECT 66.492 64.885 71.552 64.962 ;
        RECT 67.55 63.827 72.602 63.912 ;
        RECT 71.506 59.871 71.552 64.962 ;
        RECT 66.446 64.931 71.506 65.008 ;
        RECT 67.596 63.781 72.648 63.866 ;
        RECT 71.46 59.917 71.506 65.008 ;
        RECT 66.4 64.977 71.46 65.054 ;
        RECT 67.642 63.735 72.694 63.82 ;
        RECT 71.414 59.963 71.46 65.054 ;
        RECT 66.354 65.023 71.414 65.1 ;
        RECT 67.688 63.689 72.74 63.774 ;
        RECT 71.368 60.009 71.414 65.1 ;
        RECT 66.308 65.069 71.368 65.146 ;
        RECT 67.734 63.643 72.786 63.728 ;
        RECT 71.322 60.055 71.368 65.146 ;
        RECT 66.262 65.115 71.322 65.192 ;
        RECT 67.78 63.597 72.832 63.682 ;
        RECT 71.276 60.101 71.322 65.192 ;
        RECT 66.216 65.161 71.276 65.238 ;
        RECT 67.826 63.551 72.878 63.636 ;
        RECT 71.23 60.147 71.276 65.238 ;
        RECT 66.17 65.207 71.23 65.284 ;
        RECT 67.872 63.505 72.924 63.59 ;
        RECT 71.184 60.193 71.23 65.284 ;
        RECT 66.124 65.253 71.184 65.33 ;
        RECT 67.918 63.459 72.97 63.544 ;
        RECT 71.138 60.239 71.184 65.33 ;
        RECT 66.078 65.299 71.138 65.376 ;
        RECT 67.964 63.413 73.016 63.498 ;
        RECT 71.092 60.285 71.138 65.376 ;
        RECT 66.032 65.345 71.092 65.422 ;
        RECT 68.01 63.367 73.062 63.452 ;
        RECT 71.046 60.331 71.092 65.422 ;
        RECT 65.986 65.391 71.046 65.468 ;
        RECT 68.056 63.321 73.108 63.406 ;
        RECT 71 60.377 71.046 65.468 ;
        RECT 65.94 65.437 71 65.514 ;
        RECT 68.102 63.275 73.154 63.36 ;
        RECT 70.954 60.423 71 65.514 ;
        RECT 65.894 65.483 70.954 65.56 ;
        RECT 68.148 63.229 73.2 63.314 ;
        RECT 70.908 60.469 70.954 65.56 ;
        RECT 65.848 65.529 70.908 65.606 ;
        RECT 68.194 63.183 73.246 63.268 ;
        RECT 70.862 60.515 70.908 65.606 ;
        RECT 65.802 65.575 70.862 65.652 ;
        RECT 68.24 63.137 73.292 63.222 ;
        RECT 70.816 60.561 70.862 65.652 ;
        RECT 65.756 65.621 70.816 65.698 ;
        RECT 68.286 63.091 73.338 63.176 ;
        RECT 70.77 60.607 70.816 65.698 ;
        RECT 65.71 65.667 70.77 65.744 ;
        RECT 68.332 63.045 73.384 63.13 ;
        RECT 70.724 60.653 70.77 65.744 ;
        RECT 65.664 65.713 70.724 65.79 ;
        RECT 68.378 62.999 73.43 63.084 ;
        RECT 70.678 60.699 70.724 65.79 ;
        RECT 65.618 65.759 70.678 65.836 ;
        RECT 68.424 62.953 73.476 63.038 ;
        RECT 70.632 60.745 70.678 65.836 ;
        RECT 65.572 65.805 70.632 65.882 ;
        RECT 68.47 62.907 73.541 62.96 ;
        RECT 70.586 60.791 70.632 65.882 ;
        RECT 65.526 65.851 70.586 65.928 ;
        RECT 68.516 62.861 80 62.95 ;
        RECT 70.54 60.837 70.586 65.928 ;
        RECT 65.48 65.897 70.54 65.974 ;
        RECT 68.562 62.815 80 62.95 ;
        RECT 70.494 60.883 70.54 65.974 ;
        RECT 65.434 65.943 70.494 66.02 ;
        RECT 68.608 62.769 80 62.95 ;
        RECT 70.448 60.929 70.494 66.02 ;
        RECT 65.388 65.989 70.448 66.066 ;
        RECT 68.654 62.723 80 62.95 ;
        RECT 70.402 60.975 70.448 66.066 ;
        RECT 65.342 66.035 70.402 66.112 ;
        RECT 68.7 62.677 80 62.95 ;
        RECT 70.356 61.021 70.402 66.112 ;
        RECT 65.296 66.081 70.356 66.158 ;
        RECT 68.746 62.631 80 62.95 ;
        RECT 70.31 61.067 70.356 66.158 ;
        RECT 65.25 66.127 70.31 66.204 ;
        RECT 68.792 62.585 80 62.95 ;
        RECT 70.264 61.113 70.31 66.204 ;
        RECT 65.204 66.173 70.264 66.25 ;
        RECT 68.838 62.539 80 62.95 ;
        RECT 70.218 61.159 70.264 66.25 ;
        RECT 65.158 66.219 70.218 66.296 ;
        RECT 68.884 62.493 80 62.95 ;
        RECT 70.172 61.205 70.218 66.296 ;
        RECT 65.112 66.265 70.172 66.342 ;
        RECT 68.93 62.447 80 62.95 ;
        RECT 70.126 61.251 70.172 66.342 ;
        RECT 65.066 66.311 70.126 66.388 ;
        RECT 68.976 62.401 80 62.95 ;
        RECT 70.08 61.297 70.126 66.388 ;
        RECT 65.02 66.357 70.08 66.434 ;
        RECT 69.022 62.355 80 62.95 ;
        RECT 70.034 61.343 70.08 66.434 ;
        RECT 64.974 66.403 70.034 66.48 ;
        RECT 69.068 62.309 80 62.95 ;
        RECT 69.988 61.389 70.034 66.48 ;
        RECT 64.928 66.449 69.988 66.526 ;
        RECT 69.114 62.263 80 62.95 ;
        RECT 69.942 61.435 69.988 66.526 ;
        RECT 64.882 66.495 69.942 66.572 ;
        RECT 69.16 62.217 80 62.95 ;
        RECT 69.896 61.481 69.942 66.572 ;
        RECT 64.836 66.541 69.896 66.618 ;
        RECT 69.206 62.171 80 62.95 ;
        RECT 69.85 61.527 69.896 66.618 ;
        RECT 64.79 66.587 69.85 66.664 ;
        RECT 69.252 62.125 80 62.95 ;
        RECT 69.804 61.573 69.85 66.664 ;
        RECT 64.744 66.633 69.804 66.71 ;
        RECT 69.298 62.079 80 62.95 ;
        RECT 69.758 61.619 69.804 66.71 ;
        RECT 64.698 66.679 69.758 66.756 ;
        RECT 69.344 62.033 80 62.95 ;
        RECT 69.712 61.665 69.758 66.756 ;
        RECT 64.652 66.725 69.712 66.802 ;
        RECT 69.39 61.987 80 62.95 ;
        RECT 69.666 61.711 69.712 66.802 ;
        RECT 64.606 66.771 69.666 66.848 ;
        RECT 69.436 61.941 80 62.95 ;
        RECT 69.62 61.757 69.666 66.848 ;
        RECT 64.56 66.817 69.62 66.894 ;
        RECT 69.482 61.895 80 62.95 ;
        RECT 69.574 61.803 69.62 66.894 ;
        RECT 64.514 66.863 69.574 66.94 ;
        RECT 69.528 61.849 80 62.95 ;
        RECT 64.468 66.909 69.528 66.986 ;
        RECT 64.422 66.955 69.482 67.032 ;
        RECT 64.376 67.001 69.436 67.078 ;
        RECT 64.33 67.047 69.39 67.124 ;
        RECT 64.284 67.093 69.344 67.17 ;
        RECT 64.238 67.139 69.298 67.216 ;
        RECT 64.192 67.185 69.252 67.262 ;
        RECT 64.146 67.231 69.206 67.308 ;
        RECT 64.1 67.277 69.16 67.354 ;
        RECT 64.054 67.323 69.114 67.4 ;
        RECT 64.008 67.369 69.068 67.446 ;
        RECT 63.962 67.415 69.022 67.492 ;
        RECT 63.916 67.461 68.976 67.538 ;
        RECT 63.87 67.507 68.93 67.584 ;
        RECT 63.824 67.553 68.884 67.63 ;
        RECT 63.778 67.599 68.838 67.676 ;
        RECT 63.732 67.645 68.792 67.722 ;
        RECT 63.686 67.691 68.746 67.768 ;
        RECT 63.64 67.737 68.7 67.814 ;
        RECT 63.594 67.783 68.654 67.86 ;
        RECT 63.548 67.829 68.608 67.906 ;
        RECT 63.502 67.875 68.562 67.952 ;
        RECT 63.456 67.921 68.516 67.998 ;
        RECT 63.41 67.967 68.47 68.044 ;
        RECT 63.364 68.013 68.424 68.09 ;
        RECT 63.318 68.059 68.378 68.136 ;
        RECT 63.272 68.105 68.332 68.182 ;
        RECT 63.226 68.151 68.286 68.228 ;
        RECT 63.18 68.197 68.24 68.274 ;
        RECT 63.134 68.243 68.194 68.32 ;
        RECT 63.088 68.289 68.148 68.366 ;
        RECT 63.042 68.335 68.102 68.412 ;
        RECT 62.95 68.427 68.056 68.458 ;
        RECT 62.996 68.381 68.056 68.458 ;
        RECT 62.938 68.456 68.01 68.504 ;
        RECT 62.892 68.485 67.964 68.55 ;
        RECT 62.846 68.531 67.918 68.596 ;
        RECT 62.8 68.577 67.872 68.642 ;
        RECT 62.754 68.623 67.826 68.688 ;
        RECT 62.708 68.669 67.78 68.734 ;
        RECT 62.662 68.715 67.734 68.78 ;
        RECT 62.616 68.761 67.688 68.826 ;
        RECT 62.57 68.807 67.642 68.872 ;
        RECT 62.524 68.853 67.596 68.918 ;
        RECT 62.478 68.899 67.55 68.964 ;
        RECT 62.432 68.945 67.504 69.01 ;
        RECT 62.386 68.991 67.458 69.056 ;
        RECT 62.34 69.037 67.412 69.102 ;
        RECT 62.294 69.083 67.366 69.148 ;
        RECT 62.248 69.129 67.32 69.194 ;
        RECT 62.202 69.175 67.274 69.24 ;
        RECT 62.156 69.221 67.228 69.286 ;
        RECT 62.11 69.267 67.182 69.332 ;
        RECT 62.064 69.313 67.136 69.378 ;
        RECT 62.018 69.359 67.09 69.424 ;
        RECT 61.972 69.405 67.044 69.47 ;
        RECT 61.926 69.451 66.998 69.516 ;
        RECT 61.88 69.497 66.952 69.562 ;
        RECT 61.834 69.543 66.906 69.608 ;
        RECT 61.788 69.589 66.86 69.654 ;
        RECT 61.742 69.635 66.814 69.7 ;
        RECT 61.696 69.681 66.768 69.746 ;
        RECT 61.65 69.727 66.722 69.792 ;
        RECT 61.604 69.773 66.676 69.838 ;
        RECT 61.558 69.819 66.63 69.884 ;
        RECT 61.512 69.865 66.584 69.93 ;
        RECT 61.466 69.911 66.538 69.976 ;
        RECT 61.42 69.957 66.492 70.022 ;
        RECT 61.374 70.003 66.446 70.068 ;
        RECT 61.328 70.049 66.4 70.114 ;
        RECT 61.282 70.095 66.354 70.16 ;
        RECT 61.236 70.141 66.308 70.206 ;
        RECT 61.19 70.187 66.262 70.252 ;
        RECT 61.144 70.233 66.216 70.298 ;
        RECT 61.098 70.279 66.17 70.344 ;
        RECT 61.052 70.325 66.124 70.39 ;
        RECT 61.006 70.371 66.078 70.436 ;
        RECT 60.96 70.417 66.032 70.482 ;
        RECT 60.914 70.463 65.986 70.528 ;
        RECT 60.868 70.509 65.94 70.574 ;
        RECT 60.822 70.555 65.894 70.62 ;
        RECT 60.776 70.601 65.848 70.666 ;
        RECT 60.73 70.647 65.802 70.712 ;
        RECT 60.684 70.693 65.756 70.758 ;
        RECT 60.638 70.739 65.71 70.804 ;
        RECT 60.592 70.785 65.664 70.85 ;
        RECT 60.546 70.831 65.618 70.896 ;
        RECT 60.5 70.877 65.572 70.942 ;
        RECT 60.454 70.923 65.526 70.988 ;
        RECT 60.408 70.969 65.48 71.034 ;
        RECT 60.362 71.015 65.434 71.08 ;
        RECT 60.316 71.061 65.388 71.126 ;
        RECT 60.27 71.107 65.342 71.172 ;
        RECT 60.224 71.153 65.296 71.218 ;
        RECT 60.178 71.199 65.25 71.264 ;
        RECT 60.132 71.245 65.204 71.31 ;
        RECT 60.086 71.291 65.158 71.356 ;
        RECT 60.04 71.337 65.112 71.402 ;
        RECT 59.994 71.383 65.066 71.448 ;
        RECT 59.948 71.429 65.02 71.494 ;
        RECT 59.902 71.475 64.974 71.54 ;
        RECT 59.856 71.521 64.928 71.586 ;
        RECT 59.81 71.567 64.882 71.632 ;
        RECT 59.764 71.613 64.836 71.678 ;
        RECT 59.718 71.659 64.79 71.724 ;
        RECT 59.672 71.705 64.744 71.77 ;
        RECT 59.626 71.751 64.698 71.816 ;
        RECT 59.58 71.797 64.652 71.862 ;
        RECT 59.534 71.843 64.606 71.908 ;
        RECT 59.488 71.889 64.56 71.954 ;
        RECT 59.442 71.935 64.514 72 ;
        RECT 59.396 71.981 64.468 72.046 ;
        RECT 59.35 72.027 64.422 72.092 ;
        RECT 59.35 72.027 64.376 72.138 ;
        RECT 59.35 72.027 64.33 72.184 ;
        RECT 59.35 72.027 64.284 72.23 ;
        RECT 59.35 72.027 64.238 72.276 ;
        RECT 59.35 72.027 64.192 72.322 ;
        RECT 59.35 72.027 64.146 72.368 ;
        RECT 59.35 72.027 64.1 72.414 ;
        RECT 59.35 72.027 64.054 72.46 ;
        RECT 59.35 72.027 64.008 72.506 ;
        RECT 59.35 72.027 63.962 72.552 ;
        RECT 59.35 72.027 63.916 72.598 ;
        RECT 59.35 72.027 63.87 72.644 ;
        RECT 59.35 72.027 63.824 72.69 ;
        RECT 59.35 72.027 63.778 72.736 ;
        RECT 59.35 72.027 63.732 72.782 ;
        RECT 59.35 72.027 63.686 72.828 ;
        RECT 59.35 72.027 63.64 72.874 ;
        RECT 59.35 72.027 63.594 72.92 ;
        RECT 59.35 72.027 63.548 72.966 ;
        RECT 59.35 72.027 63.502 73.012 ;
        RECT 59.35 72.027 63.456 73.058 ;
        RECT 59.35 72.027 63.41 73.104 ;
        RECT 59.35 72.027 63.364 73.15 ;
        RECT 59.35 72.027 63.318 73.196 ;
        RECT 59.35 72.027 63.272 73.242 ;
        RECT 59.35 72.027 63.226 73.288 ;
        RECT 59.35 72.027 63.18 73.334 ;
        RECT 59.35 72.027 63.134 73.38 ;
        RECT 59.35 72.027 63.088 73.426 ;
        RECT 59.35 72.027 63.042 73.472 ;
        RECT 59.35 72.027 62.996 73.518 ;
        RECT 59.35 72.027 62.95 80 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 8.666 49.583 13.726 49.66 ;
        RECT 8.62 49.629 13.68 49.706 ;
        RECT 8.574 49.675 13.634 49.752 ;
        RECT 8.528 49.721 13.588 49.798 ;
        RECT 8.482 49.767 13.542 49.844 ;
        RECT 8.436 49.813 13.496 49.89 ;
        RECT 8.39 49.859 13.45 49.936 ;
        RECT 8.344 49.905 13.404 49.982 ;
        RECT 8.298 49.951 13.358 50.028 ;
        RECT 8.252 49.997 13.312 50.074 ;
        RECT 8.206 50.043 13.266 50.12 ;
        RECT 8.16 50.089 13.22 50.166 ;
        RECT 8.114 50.135 13.174 50.212 ;
        RECT 8.068 50.181 13.128 50.258 ;
        RECT 8.022 50.227 13.082 50.304 ;
        RECT 7.976 50.273 13.036 50.35 ;
        RECT 7.93 50.319 12.99 50.396 ;
        RECT 7.884 50.365 12.944 50.442 ;
        RECT 7.838 50.411 12.898 50.488 ;
        RECT 7.792 50.457 12.852 50.534 ;
        RECT 7.746 50.503 12.806 50.58 ;
        RECT 7.7 50.549 12.76 50.626 ;
        RECT 7.654 50.595 12.714 50.672 ;
        RECT 7.608 50.641 12.668 50.718 ;
        RECT 7.562 50.687 12.622 50.764 ;
        RECT 7.516 50.733 12.576 50.81 ;
        RECT 7.47 50.779 12.53 50.856 ;
        RECT 7.424 50.825 12.484 50.902 ;
        RECT 7.378 50.871 12.438 50.948 ;
        RECT 7.332 50.917 12.392 50.994 ;
        RECT 7.286 50.963 12.346 51.04 ;
        RECT 7.24 51.009 12.3 51.086 ;
        RECT 7.194 51.055 12.254 51.132 ;
        RECT 7.148 51.101 12.208 51.178 ;
        RECT 7.102 51.147 12.162 51.224 ;
        RECT 7.056 51.193 12.116 51.27 ;
        RECT 7.01 51.239 12.07 51.316 ;
        RECT 6.964 51.285 12.024 51.362 ;
        RECT 6.918 51.331 11.978 51.408 ;
        RECT 6.872 51.377 11.932 51.454 ;
        RECT 6.826 51.423 11.886 51.5 ;
        RECT 6.78 51.469 11.84 51.546 ;
        RECT 6.734 51.515 11.794 51.592 ;
        RECT 6.688 51.561 11.748 51.638 ;
        RECT 6.642 51.607 11.702 51.684 ;
        RECT 6.596 51.653 11.656 51.73 ;
        RECT 6.522 51.736 11.61 51.776 ;
        RECT 6.55 51.699 11.61 51.776 ;
        RECT 6.476 51.773 11.564 51.822 ;
        RECT 6.43 51.819 11.518 51.868 ;
        RECT 6.384 51.865 11.472 51.914 ;
        RECT 6.338 51.911 11.426 51.96 ;
        RECT 6.292 51.957 11.38 52.006 ;
        RECT 6.246 52.003 11.334 52.052 ;
        RECT 6.2 52.049 11.288 52.098 ;
        RECT 6.154 52.095 11.242 52.144 ;
        RECT 6.108 52.141 11.196 52.19 ;
        RECT 6.062 52.187 11.15 52.236 ;
        RECT 6.016 52.233 11.104 52.282 ;
        RECT 5.97 52.279 11.058 52.328 ;
        RECT 5.924 52.325 11.012 52.374 ;
        RECT 5.878 52.371 10.966 52.42 ;
        RECT 5.832 52.417 10.92 52.466 ;
        RECT 5.786 52.463 10.874 52.512 ;
        RECT 5.74 52.509 10.828 52.558 ;
        RECT 5.694 52.555 10.782 52.604 ;
        RECT 5.648 52.601 10.736 52.65 ;
        RECT 5.602 52.647 10.69 52.696 ;
        RECT 5.556 52.693 10.644 52.742 ;
        RECT 5.51 52.739 10.598 52.788 ;
        RECT 5.464 52.785 10.552 52.834 ;
        RECT 5.418 52.831 10.506 52.88 ;
        RECT 5.372 52.877 10.46 52.926 ;
        RECT 5.326 52.923 10.414 52.972 ;
        RECT 5.28 52.969 10.368 53.018 ;
        RECT 5.234 53.015 10.322 53.064 ;
        RECT 5.188 53.061 10.276 53.11 ;
        RECT 5.142 53.107 10.23 53.156 ;
        RECT 5.096 53.153 10.184 53.202 ;
        RECT 5.05 53.199 10.138 53.248 ;
        RECT 5.004 53.245 10.092 53.294 ;
        RECT 4.958 53.291 10.046 53.34 ;
        RECT 4.912 53.337 10 53.386 ;
        RECT 4.866 53.383 9.954 53.432 ;
        RECT 4.82 53.429 9.908 53.478 ;
        RECT 4.774 53.475 9.862 53.524 ;
        RECT 4.728 53.521 9.816 53.57 ;
        RECT 4.682 53.567 9.77 53.616 ;
        RECT 4.636 53.613 9.724 53.662 ;
        RECT 4.59 53.659 9.678 53.708 ;
        RECT 4.544 53.705 9.632 53.754 ;
        RECT 4.498 53.751 9.586 53.8 ;
        RECT 4.452 53.797 9.54 53.846 ;
        RECT 4.406 53.843 9.494 53.892 ;
        RECT 4.36 53.889 9.448 53.938 ;
        RECT 4.314 53.935 9.402 53.984 ;
        RECT 4.268 53.981 9.356 54.03 ;
        RECT 4.222 54.027 9.31 54.076 ;
        RECT 4.176 54.073 9.264 54.122 ;
        RECT 4.13 54.119 9.218 54.168 ;
        RECT 4.084 54.165 9.172 54.214 ;
        RECT 4.038 54.211 9.126 54.26 ;
        RECT 3.992 54.257 9.08 54.306 ;
        RECT 3.946 54.303 9.034 54.352 ;
        RECT 3.9 54.349 8.988 54.398 ;
        RECT 3.854 54.395 8.942 54.444 ;
        RECT 3.808 54.441 8.896 54.49 ;
        RECT 3.762 54.487 8.85 54.536 ;
        RECT 3.716 54.533 8.804 54.582 ;
        RECT 3.67 54.579 8.758 54.628 ;
        RECT 3.67 54.579 8.712 54.674 ;
        RECT 3.67 54.579 8.666 54.72 ;
        RECT 3.67 54.579 8.62 54.766 ;
        RECT 3.67 54.579 8.574 54.812 ;
        RECT 3.67 54.579 8.528 54.858 ;
        RECT 3.67 54.579 8.482 54.904 ;
        RECT 3.67 54.579 8.436 54.95 ;
        RECT 3.67 54.579 8.39 54.996 ;
        RECT 3.67 54.579 8.344 55.042 ;
        RECT 3.67 54.579 8.298 55.088 ;
        RECT 3.67 54.579 8.252 55.134 ;
        RECT 3.67 54.579 8.206 55.18 ;
        RECT 3.67 54.579 8.16 55.226 ;
        RECT 3.67 54.579 8.114 55.272 ;
        RECT 3.67 54.579 8.068 55.318 ;
        RECT 3.67 54.579 8.022 55.364 ;
        RECT 3.67 54.579 7.976 55.41 ;
        RECT 3.67 54.579 7.93 55.456 ;
        RECT 3.67 54.579 7.884 55.502 ;
        RECT 3.67 54.579 7.838 55.548 ;
        RECT 3.67 54.579 7.792 55.594 ;
        RECT 3.67 54.579 7.746 55.64 ;
        RECT 3.67 54.579 7.7 55.686 ;
        RECT 3.67 54.579 7.654 55.732 ;
        RECT 3.67 54.579 7.608 55.778 ;
        RECT 3.67 54.579 7.562 55.824 ;
        RECT 3.67 54.579 7.516 55.87 ;
        RECT 3.67 54.579 7.47 55.916 ;
        RECT 3.67 54.579 7.424 55.962 ;
        RECT 3.67 54.579 7.378 56.008 ;
        RECT 3.67 54.579 7.332 56.054 ;
        RECT 3.67 54.579 7.286 56.1 ;
        RECT 3.67 54.579 7.24 56.146 ;
        RECT 3.67 54.579 7.194 56.192 ;
        RECT 3.67 54.579 7.148 56.238 ;
        RECT 3.67 54.579 7.102 56.284 ;
        RECT 3.67 54.579 7.056 56.33 ;
        RECT 3.67 54.579 7.01 56.376 ;
        RECT 3.67 54.579 6.964 56.422 ;
        RECT 3.67 54.579 6.918 56.468 ;
        RECT 3.67 54.579 6.872 56.514 ;
        RECT 3.67 54.579 6.826 56.56 ;
        RECT 3.67 54.579 6.78 56.606 ;
        RECT 3.67 54.579 6.734 56.652 ;
        RECT 3.67 54.579 6.688 56.698 ;
        RECT 3.67 54.579 6.642 56.744 ;
        RECT 3.67 54.579 6.596 56.79 ;
        RECT 3.67 54.579 6.55 80 ;
        RECT 54.602 3.67 80 6.55 ;
        RECT 51.722 6.527 56.813 6.552 ;
        RECT 49.56 8.689 54.648 8.738 ;
        RECT 54.574 3.684 54.602 8.775 ;
        RECT 49.514 8.735 54.574 8.812 ;
        RECT 49.606 8.643 54.694 8.692 ;
        RECT 54.528 3.721 54.574 8.812 ;
        RECT 49.468 8.781 54.528 8.858 ;
        RECT 49.652 8.597 54.74 8.646 ;
        RECT 54.482 3.767 54.528 8.858 ;
        RECT 49.422 8.827 54.482 8.904 ;
        RECT 49.698 8.551 54.786 8.6 ;
        RECT 54.436 3.813 54.482 8.904 ;
        RECT 49.376 8.873 54.436 8.95 ;
        RECT 49.744 8.505 54.832 8.554 ;
        RECT 54.39 3.859 54.436 8.95 ;
        RECT 49.33 8.919 54.39 8.996 ;
        RECT 49.79 8.459 54.878 8.508 ;
        RECT 54.344 3.905 54.39 8.996 ;
        RECT 49.284 8.965 54.344 9.042 ;
        RECT 49.836 8.413 54.924 8.462 ;
        RECT 54.298 3.951 54.344 9.042 ;
        RECT 49.238 9.011 54.298 9.088 ;
        RECT 49.882 8.367 54.97 8.416 ;
        RECT 54.252 3.997 54.298 9.088 ;
        RECT 49.192 9.057 54.252 9.134 ;
        RECT 49.928 8.321 55.016 8.37 ;
        RECT 54.206 4.043 54.252 9.134 ;
        RECT 49.146 9.103 54.206 9.18 ;
        RECT 49.974 8.275 55.062 8.324 ;
        RECT 54.16 4.089 54.206 9.18 ;
        RECT 49.1 9.149 54.16 9.226 ;
        RECT 50.02 8.229 55.108 8.278 ;
        RECT 54.114 4.135 54.16 9.226 ;
        RECT 49.054 9.195 54.114 9.272 ;
        RECT 50.066 8.183 55.154 8.232 ;
        RECT 54.068 4.181 54.114 9.272 ;
        RECT 49.008 9.241 54.068 9.318 ;
        RECT 50.112 8.137 55.2 8.186 ;
        RECT 54.022 4.227 54.068 9.318 ;
        RECT 48.962 9.287 54.022 9.364 ;
        RECT 50.158 8.091 55.246 8.14 ;
        RECT 53.976 4.273 54.022 9.364 ;
        RECT 48.916 9.333 53.976 9.41 ;
        RECT 50.204 8.045 55.292 8.094 ;
        RECT 53.93 4.319 53.976 9.41 ;
        RECT 48.87 9.379 53.93 9.456 ;
        RECT 50.25 7.999 55.338 8.048 ;
        RECT 53.884 4.365 53.93 9.456 ;
        RECT 48.824 9.425 53.884 9.502 ;
        RECT 50.296 7.953 55.384 8.002 ;
        RECT 53.838 4.411 53.884 9.502 ;
        RECT 48.778 9.471 53.838 9.548 ;
        RECT 50.342 7.907 55.43 7.956 ;
        RECT 53.792 4.457 53.838 9.548 ;
        RECT 48.732 9.517 53.792 9.594 ;
        RECT 50.388 7.861 55.476 7.91 ;
        RECT 53.746 4.503 53.792 9.594 ;
        RECT 48.686 9.563 53.746 9.64 ;
        RECT 50.434 7.815 55.522 7.864 ;
        RECT 53.7 4.549 53.746 9.64 ;
        RECT 48.64 9.609 53.7 9.686 ;
        RECT 50.48 7.769 55.568 7.818 ;
        RECT 53.654 4.595 53.7 9.686 ;
        RECT 48.594 9.655 53.654 9.732 ;
        RECT 50.526 7.723 55.614 7.772 ;
        RECT 53.608 4.641 53.654 9.732 ;
        RECT 48.548 9.701 53.608 9.778 ;
        RECT 50.572 7.677 55.66 7.726 ;
        RECT 53.562 4.687 53.608 9.778 ;
        RECT 48.502 9.747 53.562 9.824 ;
        RECT 50.618 7.631 55.706 7.68 ;
        RECT 53.516 4.733 53.562 9.824 ;
        RECT 48.456 9.793 53.516 9.87 ;
        RECT 50.664 7.585 55.752 7.634 ;
        RECT 53.47 4.779 53.516 9.87 ;
        RECT 48.41 9.839 53.47 9.916 ;
        RECT 50.71 7.539 55.798 7.588 ;
        RECT 53.424 4.825 53.47 9.916 ;
        RECT 48.364 9.885 53.424 9.962 ;
        RECT 50.756 7.493 55.844 7.542 ;
        RECT 53.378 4.871 53.424 9.962 ;
        RECT 48.318 9.931 53.378 10.008 ;
        RECT 50.802 7.447 55.89 7.496 ;
        RECT 53.332 4.917 53.378 10.008 ;
        RECT 48.272 9.977 53.332 10.054 ;
        RECT 50.848 7.401 55.936 7.45 ;
        RECT 53.286 4.963 53.332 10.054 ;
        RECT 48.226 10.023 53.286 10.1 ;
        RECT 50.894 7.355 55.982 7.404 ;
        RECT 53.24 5.009 53.286 10.1 ;
        RECT 48.18 10.069 53.24 10.146 ;
        RECT 50.94 7.309 56.028 7.358 ;
        RECT 53.194 5.055 53.24 10.146 ;
        RECT 48.134 10.115 53.194 10.192 ;
        RECT 50.986 7.263 56.074 7.312 ;
        RECT 53.148 5.101 53.194 10.192 ;
        RECT 48.088 10.161 53.148 10.238 ;
        RECT 51.032 7.217 56.12 7.266 ;
        RECT 53.102 5.147 53.148 10.238 ;
        RECT 48.042 10.207 53.102 10.284 ;
        RECT 51.078 7.171 56.166 7.22 ;
        RECT 53.056 5.193 53.102 10.284 ;
        RECT 47.996 10.253 53.056 10.33 ;
        RECT 51.124 7.125 56.212 7.174 ;
        RECT 53.01 5.239 53.056 10.33 ;
        RECT 47.95 10.299 53.01 10.376 ;
        RECT 51.17 7.079 56.258 7.128 ;
        RECT 52.964 5.285 53.01 10.376 ;
        RECT 47.904 10.345 52.964 10.422 ;
        RECT 51.216 7.033 56.304 7.082 ;
        RECT 52.918 5.331 52.964 10.422 ;
        RECT 47.858 10.391 52.918 10.468 ;
        RECT 51.262 6.987 56.35 7.036 ;
        RECT 52.872 5.377 52.918 10.468 ;
        RECT 47.812 10.437 52.872 10.514 ;
        RECT 51.308 6.941 56.396 6.99 ;
        RECT 52.826 5.423 52.872 10.514 ;
        RECT 47.766 10.483 52.826 10.56 ;
        RECT 51.354 6.895 56.442 6.944 ;
        RECT 52.78 5.469 52.826 10.56 ;
        RECT 47.72 10.529 52.78 10.606 ;
        RECT 51.4 6.849 56.488 6.898 ;
        RECT 52.734 5.515 52.78 10.606 ;
        RECT 47.674 10.575 52.734 10.652 ;
        RECT 51.446 6.803 56.534 6.852 ;
        RECT 52.688 5.561 52.734 10.652 ;
        RECT 47.628 10.621 52.688 10.698 ;
        RECT 51.492 6.757 56.58 6.806 ;
        RECT 52.642 5.607 52.688 10.698 ;
        RECT 47.582 10.667 52.642 10.744 ;
        RECT 51.538 6.711 56.626 6.76 ;
        RECT 52.596 5.653 52.642 10.744 ;
        RECT 47.536 10.713 52.596 10.79 ;
        RECT 51.584 6.665 56.672 6.714 ;
        RECT 52.55 5.699 52.596 10.79 ;
        RECT 47.49 10.759 52.55 10.836 ;
        RECT 51.63 6.619 56.718 6.668 ;
        RECT 52.504 5.745 52.55 10.836 ;
        RECT 47.444 10.805 52.504 10.882 ;
        RECT 51.676 6.573 56.764 6.622 ;
        RECT 52.458 5.791 52.504 10.882 ;
        RECT 47.398 10.851 52.458 10.928 ;
        RECT 51.722 6.527 56.81 6.576 ;
        RECT 52.412 5.837 52.458 10.928 ;
        RECT 47.352 10.897 52.412 10.974 ;
        RECT 51.768 6.481 80 6.55 ;
        RECT 52.366 5.883 52.412 10.974 ;
        RECT 47.306 10.943 52.366 11.02 ;
        RECT 51.814 6.435 80 6.55 ;
        RECT 52.32 5.929 52.366 11.02 ;
        RECT 47.26 10.989 52.32 11.066 ;
        RECT 51.86 6.389 80 6.55 ;
        RECT 52.274 5.975 52.32 11.066 ;
        RECT 47.214 11.035 52.274 11.112 ;
        RECT 51.906 6.343 80 6.55 ;
        RECT 52.228 6.021 52.274 11.112 ;
        RECT 47.168 11.081 52.228 11.158 ;
        RECT 51.952 6.297 80 6.55 ;
        RECT 52.182 6.067 52.228 11.158 ;
        RECT 47.122 11.127 52.182 11.204 ;
        RECT 51.998 6.251 80 6.55 ;
        RECT 52.136 6.113 52.182 11.204 ;
        RECT 47.076 11.173 52.136 11.25 ;
        RECT 52.044 6.205 80 6.55 ;
        RECT 52.09 6.159 52.136 11.25 ;
        RECT 47.03 11.219 52.09 11.296 ;
        RECT 46.984 11.265 52.044 11.342 ;
        RECT 46.938 11.311 51.998 11.388 ;
        RECT 46.892 11.357 51.952 11.434 ;
        RECT 46.846 11.403 51.906 11.48 ;
        RECT 46.8 11.449 51.86 11.526 ;
        RECT 46.754 11.495 51.814 11.572 ;
        RECT 46.708 11.541 51.768 11.618 ;
        RECT 46.662 11.587 51.722 11.664 ;
        RECT 46.616 11.633 51.676 11.71 ;
        RECT 46.57 11.679 51.63 11.756 ;
        RECT 46.524 11.725 51.584 11.802 ;
        RECT 46.478 11.771 51.538 11.848 ;
        RECT 46.432 11.817 51.492 11.894 ;
        RECT 46.386 11.863 51.446 11.94 ;
        RECT 46.34 11.909 51.4 11.986 ;
        RECT 46.294 11.955 51.354 12.032 ;
        RECT 46.248 12.001 51.308 12.078 ;
        RECT 46.202 12.047 51.262 12.124 ;
        RECT 46.156 12.093 51.216 12.17 ;
        RECT 46.11 12.139 51.17 12.216 ;
        RECT 46.064 12.185 51.124 12.262 ;
        RECT 46.018 12.231 51.078 12.308 ;
        RECT 45.972 12.277 51.032 12.354 ;
        RECT 45.926 12.323 50.986 12.4 ;
        RECT 45.88 12.369 50.94 12.446 ;
        RECT 45.834 12.415 50.894 12.492 ;
        RECT 45.788 12.461 50.848 12.538 ;
        RECT 45.742 12.507 50.802 12.584 ;
        RECT 45.696 12.553 50.756 12.63 ;
        RECT 45.65 12.599 50.71 12.676 ;
        RECT 45.604 12.645 50.664 12.722 ;
        RECT 45.558 12.691 50.618 12.768 ;
        RECT 45.512 12.737 50.572 12.814 ;
        RECT 45.466 12.783 50.526 12.86 ;
        RECT 45.42 12.829 50.48 12.906 ;
        RECT 45.374 12.875 50.434 12.952 ;
        RECT 45.328 12.921 50.388 12.998 ;
        RECT 45.282 12.967 50.342 13.044 ;
        RECT 45.236 13.013 50.296 13.09 ;
        RECT 45.19 13.059 50.25 13.136 ;
        RECT 45.144 13.105 50.204 13.182 ;
        RECT 45.098 13.151 50.158 13.228 ;
        RECT 45.052 13.197 50.112 13.274 ;
        RECT 45.006 13.243 50.066 13.32 ;
        RECT 44.96 13.289 50.02 13.366 ;
        RECT 44.914 13.335 49.974 13.412 ;
        RECT 44.868 13.381 49.928 13.458 ;
        RECT 44.822 13.427 49.882 13.504 ;
        RECT 44.776 13.473 49.836 13.55 ;
        RECT 44.73 13.519 49.79 13.596 ;
        RECT 44.684 13.565 49.744 13.642 ;
        RECT 44.638 13.611 49.698 13.688 ;
        RECT 44.592 13.657 49.652 13.734 ;
        RECT 44.546 13.703 49.606 13.78 ;
        RECT 44.5 13.749 49.56 13.826 ;
        RECT 44.454 13.795 49.514 13.872 ;
        RECT 44.408 13.841 49.468 13.918 ;
        RECT 44.362 13.887 49.422 13.964 ;
        RECT 44.316 13.933 49.376 14.01 ;
        RECT 44.27 13.979 49.33 14.056 ;
        RECT 44.224 14.025 49.284 14.102 ;
        RECT 44.178 14.071 49.238 14.148 ;
        RECT 44.132 14.117 49.192 14.194 ;
        RECT 44.086 14.163 49.146 14.24 ;
        RECT 44.04 14.209 49.1 14.286 ;
        RECT 43.994 14.255 49.054 14.332 ;
        RECT 43.948 14.301 49.008 14.378 ;
        RECT 43.902 14.347 48.962 14.424 ;
        RECT 43.856 14.393 48.916 14.47 ;
        RECT 43.81 14.439 48.87 14.516 ;
        RECT 43.764 14.485 48.824 14.562 ;
        RECT 43.718 14.531 48.778 14.608 ;
        RECT 43.672 14.577 48.732 14.654 ;
        RECT 43.626 14.623 48.686 14.7 ;
        RECT 43.58 14.669 48.64 14.746 ;
        RECT 43.534 14.715 48.594 14.792 ;
        RECT 43.488 14.761 48.548 14.838 ;
        RECT 43.442 14.807 48.502 14.884 ;
        RECT 43.396 14.853 48.456 14.93 ;
        RECT 43.35 14.899 48.41 14.976 ;
        RECT 43.304 14.945 48.364 15.022 ;
        RECT 43.258 14.991 48.318 15.068 ;
        RECT 43.212 15.037 48.272 15.114 ;
        RECT 43.166 15.083 48.226 15.16 ;
        RECT 43.12 15.129 48.18 15.206 ;
        RECT 43.074 15.175 48.134 15.252 ;
        RECT 43.028 15.221 48.088 15.298 ;
        RECT 42.982 15.267 48.042 15.344 ;
        RECT 42.936 15.313 47.996 15.39 ;
        RECT 42.89 15.359 47.95 15.436 ;
        RECT 42.844 15.405 47.904 15.482 ;
        RECT 42.798 15.451 47.858 15.528 ;
        RECT 42.752 15.497 47.812 15.574 ;
        RECT 42.706 15.543 47.766 15.62 ;
        RECT 42.66 15.589 47.72 15.666 ;
        RECT 42.614 15.635 47.674 15.712 ;
        RECT 42.568 15.681 47.628 15.758 ;
        RECT 42.522 15.727 47.582 15.804 ;
        RECT 42.476 15.773 47.536 15.85 ;
        RECT 42.43 15.819 47.49 15.896 ;
        RECT 42.384 15.865 47.444 15.942 ;
        RECT 42.338 15.911 47.398 15.988 ;
        RECT 42.292 15.957 47.352 16.034 ;
        RECT 42.246 16.003 47.306 16.08 ;
        RECT 42.2 16.049 47.26 16.126 ;
        RECT 42.154 16.095 47.214 16.172 ;
        RECT 42.108 16.141 47.168 16.218 ;
        RECT 42.062 16.187 47.122 16.264 ;
        RECT 42.016 16.233 47.076 16.31 ;
        RECT 41.97 16.279 47.03 16.356 ;
        RECT 41.924 16.325 46.984 16.402 ;
        RECT 41.878 16.371 46.938 16.448 ;
        RECT 41.832 16.417 46.892 16.494 ;
        RECT 41.786 16.463 46.846 16.54 ;
        RECT 41.74 16.509 46.8 16.586 ;
        RECT 41.694 16.555 46.754 16.632 ;
        RECT 41.648 16.601 46.708 16.678 ;
        RECT 41.602 16.647 46.662 16.724 ;
        RECT 41.556 16.693 46.616 16.77 ;
        RECT 41.51 16.739 46.57 16.816 ;
        RECT 41.464 16.785 46.524 16.862 ;
        RECT 41.418 16.831 46.478 16.908 ;
        RECT 41.372 16.877 46.432 16.954 ;
        RECT 41.326 16.923 46.386 17 ;
        RECT 41.28 16.969 46.34 17.046 ;
        RECT 41.234 17.015 46.294 17.092 ;
        RECT 41.188 17.061 46.248 17.138 ;
        RECT 41.142 17.107 46.202 17.184 ;
        RECT 41.096 17.153 46.156 17.23 ;
        RECT 41.05 17.199 46.11 17.276 ;
        RECT 41.004 17.245 46.064 17.322 ;
        RECT 40.958 17.291 46.018 17.368 ;
        RECT 40.912 17.337 45.972 17.414 ;
        RECT 40.866 17.383 45.926 17.46 ;
        RECT 40.82 17.429 45.88 17.506 ;
        RECT 40.774 17.475 45.834 17.552 ;
        RECT 40.728 17.521 45.788 17.598 ;
        RECT 40.682 17.567 45.742 17.644 ;
        RECT 40.636 17.613 45.696 17.69 ;
        RECT 40.59 17.659 45.65 17.736 ;
        RECT 40.544 17.705 45.604 17.782 ;
        RECT 40.498 17.751 45.558 17.828 ;
        RECT 40.452 17.797 45.512 17.874 ;
        RECT 40.406 17.843 45.466 17.92 ;
        RECT 40.36 17.889 45.42 17.966 ;
        RECT 40.314 17.935 45.374 18.012 ;
        RECT 40.268 17.981 45.328 18.058 ;
        RECT 40.222 18.027 45.282 18.104 ;
        RECT 40.176 18.073 45.236 18.15 ;
        RECT 40.13 18.119 45.19 18.196 ;
        RECT 40.084 18.165 45.144 18.242 ;
        RECT 40.038 18.211 45.098 18.288 ;
        RECT 39.992 18.257 45.052 18.334 ;
        RECT 39.946 18.303 45.006 18.38 ;
        RECT 39.9 18.349 44.96 18.426 ;
        RECT 39.854 18.395 44.914 18.472 ;
        RECT 39.808 18.441 44.868 18.518 ;
        RECT 39.762 18.487 44.822 18.564 ;
        RECT 39.716 18.533 44.776 18.61 ;
        RECT 39.67 18.579 44.73 18.656 ;
        RECT 39.624 18.625 44.684 18.702 ;
        RECT 39.578 18.671 44.638 18.748 ;
        RECT 39.532 18.717 44.592 18.794 ;
        RECT 39.486 18.763 44.546 18.84 ;
        RECT 39.44 18.809 44.5 18.886 ;
        RECT 39.394 18.855 44.454 18.932 ;
        RECT 39.348 18.901 44.408 18.978 ;
        RECT 39.302 18.947 44.362 19.024 ;
        RECT 39.256 18.993 44.316 19.07 ;
        RECT 39.21 19.039 44.27 19.116 ;
        RECT 39.164 19.085 44.224 19.162 ;
        RECT 39.118 19.131 44.178 19.208 ;
        RECT 39.072 19.177 44.132 19.254 ;
        RECT 39.026 19.223 44.086 19.3 ;
        RECT 38.98 19.269 44.04 19.346 ;
        RECT 38.934 19.315 43.994 19.392 ;
        RECT 38.888 19.361 43.948 19.438 ;
        RECT 38.842 19.407 43.902 19.484 ;
        RECT 38.796 19.453 43.856 19.53 ;
        RECT 38.75 19.499 43.81 19.576 ;
        RECT 38.704 19.545 43.764 19.622 ;
        RECT 38.658 19.591 43.718 19.668 ;
        RECT 38.612 19.637 43.672 19.714 ;
        RECT 38.566 19.683 43.626 19.76 ;
        RECT 38.52 19.729 43.58 19.806 ;
        RECT 38.474 19.775 43.534 19.852 ;
        RECT 38.428 19.821 43.488 19.898 ;
        RECT 38.382 19.867 43.442 19.944 ;
        RECT 38.336 19.913 43.396 19.99 ;
        RECT 38.29 19.959 43.35 20.036 ;
        RECT 38.244 20.005 43.304 20.082 ;
        RECT 38.198 20.051 43.258 20.128 ;
        RECT 38.152 20.097 43.212 20.174 ;
        RECT 38.106 20.143 43.166 20.22 ;
        RECT 38.06 20.189 43.12 20.266 ;
        RECT 38.014 20.235 43.074 20.312 ;
        RECT 37.968 20.281 43.028 20.358 ;
        RECT 37.922 20.327 42.982 20.404 ;
        RECT 37.876 20.373 42.936 20.45 ;
        RECT 37.83 20.419 42.89 20.496 ;
        RECT 37.784 20.465 42.844 20.542 ;
        RECT 37.738 20.511 42.798 20.588 ;
        RECT 37.692 20.557 42.752 20.634 ;
        RECT 37.646 20.603 42.706 20.68 ;
        RECT 37.6 20.649 42.66 20.726 ;
        RECT 37.554 20.695 42.614 20.772 ;
        RECT 37.508 20.741 42.568 20.818 ;
        RECT 37.462 20.787 42.522 20.864 ;
        RECT 37.416 20.833 42.476 20.91 ;
        RECT 37.37 20.879 42.43 20.956 ;
        RECT 37.324 20.925 42.384 21.002 ;
        RECT 37.278 20.971 42.338 21.048 ;
        RECT 37.232 21.017 42.292 21.094 ;
        RECT 37.186 21.063 42.246 21.14 ;
        RECT 37.14 21.109 42.2 21.186 ;
        RECT 37.094 21.155 42.154 21.232 ;
        RECT 37.048 21.201 42.108 21.278 ;
        RECT 37.002 21.247 42.062 21.324 ;
        RECT 36.956 21.293 42.016 21.37 ;
        RECT 36.91 21.339 41.97 21.416 ;
        RECT 36.864 21.385 41.924 21.462 ;
        RECT 36.818 21.431 41.878 21.508 ;
        RECT 36.772 21.477 41.832 21.554 ;
        RECT 36.726 21.523 41.786 21.6 ;
        RECT 36.68 21.569 41.74 21.646 ;
        RECT 36.634 21.615 41.694 21.692 ;
        RECT 36.588 21.661 41.648 21.738 ;
        RECT 36.542 21.707 41.602 21.784 ;
        RECT 36.496 21.753 41.556 21.83 ;
        RECT 36.45 21.799 41.51 21.876 ;
        RECT 36.404 21.845 41.464 21.922 ;
        RECT 36.358 21.891 41.418 21.968 ;
        RECT 36.312 21.937 41.372 22.014 ;
        RECT 36.266 21.983 41.326 22.06 ;
        RECT 36.22 22.029 41.28 22.106 ;
        RECT 36.174 22.075 41.234 22.152 ;
        RECT 36.128 22.121 41.188 22.198 ;
        RECT 36.082 22.167 41.142 22.244 ;
        RECT 36.036 22.213 41.096 22.29 ;
        RECT 35.99 22.259 41.05 22.336 ;
        RECT 35.944 22.305 41.004 22.382 ;
        RECT 35.898 22.351 40.958 22.428 ;
        RECT 35.852 22.397 40.912 22.474 ;
        RECT 35.806 22.443 40.866 22.52 ;
        RECT 35.76 22.489 40.82 22.566 ;
        RECT 35.714 22.535 40.774 22.612 ;
        RECT 35.668 22.581 40.728 22.658 ;
        RECT 35.622 22.627 40.682 22.704 ;
        RECT 35.576 22.673 40.636 22.75 ;
        RECT 35.53 22.719 40.59 22.796 ;
        RECT 35.484 22.765 40.544 22.842 ;
        RECT 35.438 22.811 40.498 22.888 ;
        RECT 35.392 22.857 40.452 22.934 ;
        RECT 35.346 22.903 40.406 22.98 ;
        RECT 35.3 22.949 40.36 23.026 ;
        RECT 35.254 22.995 40.314 23.072 ;
        RECT 35.208 23.041 40.268 23.118 ;
        RECT 35.162 23.087 40.222 23.164 ;
        RECT 35.116 23.133 40.176 23.21 ;
        RECT 35.07 23.179 40.13 23.256 ;
        RECT 35.024 23.225 40.084 23.302 ;
        RECT 34.978 23.271 40.038 23.348 ;
        RECT 34.932 23.317 39.992 23.394 ;
        RECT 34.886 23.363 39.946 23.44 ;
        RECT 34.84 23.409 39.9 23.486 ;
        RECT 34.794 23.455 39.854 23.532 ;
        RECT 34.748 23.501 39.808 23.578 ;
        RECT 34.702 23.547 39.762 23.624 ;
        RECT 34.656 23.593 39.716 23.67 ;
        RECT 34.61 23.639 39.67 23.716 ;
        RECT 34.564 23.685 39.624 23.762 ;
        RECT 34.518 23.731 39.578 23.808 ;
        RECT 34.472 23.777 39.532 23.854 ;
        RECT 34.426 23.823 39.486 23.9 ;
        RECT 34.38 23.869 39.44 23.946 ;
        RECT 34.334 23.915 39.394 23.992 ;
        RECT 34.288 23.961 39.348 24.038 ;
        RECT 34.242 24.007 39.302 24.084 ;
        RECT 34.196 24.053 39.256 24.13 ;
        RECT 34.15 24.099 39.21 24.176 ;
        RECT 34.104 24.145 39.164 24.222 ;
        RECT 34.058 24.191 39.118 24.268 ;
        RECT 34.012 24.237 39.072 24.314 ;
        RECT 33.966 24.283 39.026 24.36 ;
        RECT 33.92 24.329 38.98 24.406 ;
        RECT 33.874 24.375 38.934 24.452 ;
        RECT 33.828 24.421 38.888 24.498 ;
        RECT 33.782 24.467 38.842 24.544 ;
        RECT 33.736 24.513 38.796 24.59 ;
        RECT 33.69 24.559 38.75 24.636 ;
        RECT 33.644 24.605 38.704 24.682 ;
        RECT 33.598 24.651 38.658 24.728 ;
        RECT 33.552 24.697 38.612 24.774 ;
        RECT 33.506 24.743 38.566 24.82 ;
        RECT 33.46 24.789 38.52 24.866 ;
        RECT 33.414 24.835 38.474 24.912 ;
        RECT 33.368 24.881 38.428 24.958 ;
        RECT 33.322 24.927 38.382 25.004 ;
        RECT 33.276 24.973 38.336 25.05 ;
        RECT 33.23 25.019 38.29 25.096 ;
        RECT 33.184 25.065 38.244 25.142 ;
        RECT 33.138 25.111 38.198 25.188 ;
        RECT 33.092 25.157 38.152 25.234 ;
        RECT 33.046 25.203 38.106 25.28 ;
        RECT 33 25.249 38.06 25.326 ;
        RECT 32.954 25.295 38.014 25.372 ;
        RECT 32.908 25.341 37.968 25.418 ;
        RECT 32.862 25.387 37.922 25.464 ;
        RECT 32.816 25.433 37.876 25.51 ;
        RECT 32.77 25.479 37.83 25.556 ;
        RECT 32.724 25.525 37.784 25.602 ;
        RECT 32.678 25.571 37.738 25.648 ;
        RECT 32.632 25.617 37.692 25.694 ;
        RECT 32.586 25.663 37.646 25.74 ;
        RECT 32.54 25.709 37.6 25.786 ;
        RECT 32.494 25.755 37.554 25.832 ;
        RECT 32.448 25.801 37.508 25.878 ;
        RECT 32.402 25.847 37.462 25.924 ;
        RECT 32.356 25.893 37.416 25.97 ;
        RECT 32.31 25.939 37.37 26.016 ;
        RECT 32.264 25.985 37.324 26.062 ;
        RECT 32.218 26.031 37.278 26.108 ;
        RECT 32.172 26.077 37.232 26.154 ;
        RECT 32.126 26.123 37.186 26.2 ;
        RECT 32.08 26.169 37.14 26.246 ;
        RECT 32.034 26.215 37.094 26.292 ;
        RECT 31.988 26.261 37.048 26.338 ;
        RECT 31.942 26.307 37.002 26.384 ;
        RECT 31.896 26.353 36.956 26.43 ;
        RECT 31.85 26.399 36.91 26.476 ;
        RECT 31.804 26.445 36.864 26.522 ;
        RECT 31.758 26.491 36.818 26.568 ;
        RECT 31.712 26.537 36.772 26.614 ;
        RECT 31.666 26.583 36.726 26.66 ;
        RECT 31.62 26.629 36.68 26.706 ;
        RECT 31.574 26.675 36.634 26.752 ;
        RECT 31.528 26.721 36.588 26.798 ;
        RECT 31.482 26.767 36.542 26.844 ;
        RECT 31.436 26.813 36.496 26.89 ;
        RECT 31.39 26.859 36.45 26.936 ;
        RECT 31.344 26.905 36.404 26.982 ;
        RECT 31.298 26.951 36.358 27.028 ;
        RECT 31.252 26.997 36.312 27.074 ;
        RECT 31.206 27.043 36.266 27.12 ;
        RECT 31.16 27.089 36.22 27.166 ;
        RECT 31.114 27.135 36.174 27.212 ;
        RECT 31.068 27.181 36.128 27.258 ;
        RECT 31.022 27.227 36.082 27.304 ;
        RECT 30.976 27.273 36.036 27.35 ;
        RECT 30.93 27.319 35.99 27.396 ;
        RECT 30.884 27.365 35.944 27.442 ;
        RECT 30.838 27.411 35.898 27.488 ;
        RECT 30.792 27.457 35.852 27.534 ;
        RECT 30.746 27.503 35.806 27.58 ;
        RECT 30.7 27.549 35.76 27.626 ;
        RECT 30.654 27.595 35.714 27.672 ;
        RECT 30.608 27.641 35.668 27.718 ;
        RECT 30.562 27.687 35.622 27.764 ;
        RECT 30.516 27.733 35.576 27.81 ;
        RECT 30.47 27.779 35.53 27.856 ;
        RECT 30.424 27.825 35.484 27.902 ;
        RECT 30.378 27.871 35.438 27.948 ;
        RECT 30.332 27.917 35.392 27.994 ;
        RECT 30.286 27.963 35.346 28.04 ;
        RECT 30.24 28.009 35.3 28.086 ;
        RECT 30.194 28.055 35.254 28.132 ;
        RECT 30.148 28.101 35.208 28.178 ;
        RECT 30.102 28.147 35.162 28.224 ;
        RECT 30.056 28.193 35.116 28.27 ;
        RECT 30.01 28.239 35.07 28.316 ;
        RECT 29.964 28.285 35.024 28.362 ;
        RECT 29.918 28.331 34.978 28.408 ;
        RECT 29.872 28.377 34.932 28.454 ;
        RECT 29.826 28.423 34.886 28.5 ;
        RECT 29.78 28.469 34.84 28.546 ;
        RECT 29.734 28.515 34.794 28.592 ;
        RECT 29.688 28.561 34.748 28.638 ;
        RECT 29.642 28.607 34.702 28.684 ;
        RECT 29.596 28.653 34.656 28.73 ;
        RECT 29.55 28.699 34.61 28.776 ;
        RECT 29.504 28.745 34.564 28.822 ;
        RECT 29.458 28.791 34.518 28.868 ;
        RECT 29.412 28.837 34.472 28.914 ;
        RECT 29.366 28.883 34.426 28.96 ;
        RECT 29.32 28.929 34.38 29.006 ;
        RECT 29.274 28.975 34.334 29.052 ;
        RECT 29.228 29.021 34.288 29.098 ;
        RECT 29.182 29.067 34.242 29.144 ;
        RECT 29.136 29.113 34.196 29.19 ;
        RECT 29.09 29.159 34.15 29.236 ;
        RECT 29.044 29.205 34.104 29.282 ;
        RECT 28.998 29.251 34.058 29.328 ;
        RECT 28.952 29.297 34.012 29.374 ;
        RECT 28.906 29.343 33.966 29.42 ;
        RECT 28.86 29.389 33.92 29.466 ;
        RECT 28.814 29.435 33.874 29.512 ;
        RECT 28.768 29.481 33.828 29.558 ;
        RECT 28.722 29.527 33.782 29.604 ;
        RECT 28.676 29.573 33.736 29.65 ;
        RECT 28.63 29.619 33.69 29.696 ;
        RECT 28.584 29.665 33.644 29.742 ;
        RECT 28.538 29.711 33.598 29.788 ;
        RECT 28.492 29.757 33.552 29.834 ;
        RECT 28.446 29.803 33.506 29.88 ;
        RECT 28.4 29.849 33.46 29.926 ;
        RECT 28.354 29.895 33.414 29.972 ;
        RECT 28.308 29.941 33.368 30.018 ;
        RECT 28.262 29.987 33.322 30.064 ;
        RECT 28.216 30.033 33.276 30.11 ;
        RECT 28.17 30.079 33.23 30.156 ;
        RECT 28.124 30.125 33.184 30.202 ;
        RECT 28.078 30.171 33.138 30.248 ;
        RECT 28.032 30.217 33.092 30.294 ;
        RECT 27.986 30.263 33.046 30.34 ;
        RECT 27.94 30.309 33 30.386 ;
        RECT 27.894 30.355 32.954 30.432 ;
        RECT 27.848 30.401 32.908 30.478 ;
        RECT 27.802 30.447 32.862 30.524 ;
        RECT 27.756 30.493 32.816 30.57 ;
        RECT 27.71 30.539 32.77 30.616 ;
        RECT 27.664 30.585 32.724 30.662 ;
        RECT 27.618 30.631 32.678 30.708 ;
        RECT 27.572 30.677 32.632 30.754 ;
        RECT 27.526 30.723 32.586 30.8 ;
        RECT 27.48 30.769 32.54 30.846 ;
        RECT 27.434 30.815 32.494 30.892 ;
        RECT 27.388 30.861 32.448 30.938 ;
        RECT 27.342 30.907 32.402 30.984 ;
        RECT 27.296 30.953 32.356 31.03 ;
        RECT 27.25 30.999 32.31 31.076 ;
        RECT 27.204 31.045 32.264 31.122 ;
        RECT 27.158 31.091 32.218 31.168 ;
        RECT 27.112 31.137 32.172 31.214 ;
        RECT 27.066 31.183 32.126 31.26 ;
        RECT 27.02 31.229 32.08 31.306 ;
        RECT 26.974 31.275 32.034 31.352 ;
        RECT 26.928 31.321 31.988 31.398 ;
        RECT 26.882 31.367 31.942 31.444 ;
        RECT 26.836 31.413 31.896 31.49 ;
        RECT 26.79 31.459 31.85 31.536 ;
        RECT 26.744 31.505 31.804 31.582 ;
        RECT 26.698 31.551 31.758 31.628 ;
        RECT 26.652 31.597 31.712 31.674 ;
        RECT 26.606 31.643 31.666 31.72 ;
        RECT 26.56 31.689 31.62 31.766 ;
        RECT 26.514 31.735 31.574 31.812 ;
        RECT 26.468 31.781 31.528 31.858 ;
        RECT 26.422 31.827 31.482 31.904 ;
        RECT 26.376 31.873 31.436 31.95 ;
        RECT 26.33 31.919 31.39 31.996 ;
        RECT 26.284 31.965 31.344 32.042 ;
        RECT 26.238 32.011 31.298 32.088 ;
        RECT 26.192 32.057 31.252 32.134 ;
        RECT 26.146 32.103 31.206 32.18 ;
        RECT 26.1 32.149 31.16 32.226 ;
        RECT 26.054 32.195 31.114 32.272 ;
        RECT 26.008 32.241 31.068 32.318 ;
        RECT 25.962 32.287 31.022 32.364 ;
        RECT 25.916 32.333 30.976 32.41 ;
        RECT 25.87 32.379 30.93 32.456 ;
        RECT 25.824 32.425 30.884 32.502 ;
        RECT 25.778 32.471 30.838 32.548 ;
        RECT 25.732 32.517 30.792 32.594 ;
        RECT 25.686 32.563 30.746 32.64 ;
        RECT 25.64 32.609 30.7 32.686 ;
        RECT 25.594 32.655 30.654 32.732 ;
        RECT 25.548 32.701 30.608 32.778 ;
        RECT 25.502 32.747 30.562 32.824 ;
        RECT 25.456 32.793 30.516 32.87 ;
        RECT 25.41 32.839 30.47 32.916 ;
        RECT 25.364 32.885 30.424 32.962 ;
        RECT 25.318 32.931 30.378 33.008 ;
        RECT 25.272 32.977 30.332 33.054 ;
        RECT 25.226 33.023 30.286 33.1 ;
        RECT 25.18 33.069 30.24 33.146 ;
        RECT 25.134 33.115 30.194 33.192 ;
        RECT 25.088 33.161 30.148 33.238 ;
        RECT 25.042 33.207 30.102 33.284 ;
        RECT 24.996 33.253 30.056 33.33 ;
        RECT 24.95 33.299 30.01 33.376 ;
        RECT 24.904 33.345 29.964 33.422 ;
        RECT 24.858 33.391 29.918 33.468 ;
        RECT 24.812 33.437 29.872 33.514 ;
        RECT 24.766 33.483 29.826 33.56 ;
        RECT 24.72 33.529 29.78 33.606 ;
        RECT 24.674 33.575 29.734 33.652 ;
        RECT 24.628 33.621 29.688 33.698 ;
        RECT 24.582 33.667 29.642 33.744 ;
        RECT 24.536 33.713 29.596 33.79 ;
        RECT 24.49 33.759 29.55 33.836 ;
        RECT 24.444 33.805 29.504 33.882 ;
        RECT 24.398 33.851 29.458 33.928 ;
        RECT 24.352 33.897 29.412 33.974 ;
        RECT 24.306 33.943 29.366 34.02 ;
        RECT 24.26 33.989 29.32 34.066 ;
        RECT 24.214 34.035 29.274 34.112 ;
        RECT 24.168 34.081 29.228 34.158 ;
        RECT 24.122 34.127 29.182 34.204 ;
        RECT 24.076 34.173 29.136 34.25 ;
        RECT 24.03 34.219 29.09 34.296 ;
        RECT 23.984 34.265 29.044 34.342 ;
        RECT 23.938 34.311 28.998 34.388 ;
        RECT 23.892 34.357 28.952 34.434 ;
        RECT 23.846 34.403 28.906 34.48 ;
        RECT 23.8 34.449 28.86 34.526 ;
        RECT 23.754 34.495 28.814 34.572 ;
        RECT 23.708 34.541 28.768 34.618 ;
        RECT 23.662 34.587 28.722 34.664 ;
        RECT 23.616 34.633 28.676 34.71 ;
        RECT 23.57 34.679 28.63 34.756 ;
        RECT 23.524 34.725 28.584 34.802 ;
        RECT 23.478 34.771 28.538 34.848 ;
        RECT 23.432 34.817 28.492 34.894 ;
        RECT 23.386 34.863 28.446 34.94 ;
        RECT 23.34 34.909 28.4 34.986 ;
        RECT 23.294 34.955 28.354 35.032 ;
        RECT 23.248 35.001 28.308 35.078 ;
        RECT 23.202 35.047 28.262 35.124 ;
        RECT 23.156 35.093 28.216 35.17 ;
        RECT 23.11 35.139 28.17 35.216 ;
        RECT 23.064 35.185 28.124 35.262 ;
        RECT 23.018 35.231 28.078 35.308 ;
        RECT 22.972 35.277 28.032 35.354 ;
        RECT 22.926 35.323 27.986 35.4 ;
        RECT 22.88 35.369 27.94 35.446 ;
        RECT 22.834 35.415 27.894 35.492 ;
        RECT 22.788 35.461 27.848 35.538 ;
        RECT 22.742 35.507 27.802 35.584 ;
        RECT 22.696 35.553 27.756 35.63 ;
        RECT 22.65 35.599 27.71 35.676 ;
        RECT 22.604 35.645 27.664 35.722 ;
        RECT 22.558 35.691 27.618 35.768 ;
        RECT 22.512 35.737 27.572 35.814 ;
        RECT 22.466 35.783 27.526 35.86 ;
        RECT 22.42 35.829 27.48 35.906 ;
        RECT 22.374 35.875 27.434 35.952 ;
        RECT 22.328 35.921 27.388 35.998 ;
        RECT 22.282 35.967 27.342 36.044 ;
        RECT 22.236 36.013 27.296 36.09 ;
        RECT 22.19 36.059 27.25 36.136 ;
        RECT 22.144 36.105 27.204 36.182 ;
        RECT 22.098 36.151 27.158 36.228 ;
        RECT 22.052 36.197 27.112 36.274 ;
        RECT 22.006 36.243 27.066 36.32 ;
        RECT 21.96 36.289 27.02 36.366 ;
        RECT 21.914 36.335 26.974 36.412 ;
        RECT 21.868 36.381 26.928 36.458 ;
        RECT 21.822 36.427 26.882 36.504 ;
        RECT 21.776 36.473 26.836 36.55 ;
        RECT 21.73 36.519 26.79 36.596 ;
        RECT 21.684 36.565 26.744 36.642 ;
        RECT 21.638 36.611 26.698 36.688 ;
        RECT 21.592 36.657 26.652 36.734 ;
        RECT 21.546 36.703 26.606 36.78 ;
        RECT 21.5 36.749 26.56 36.826 ;
        RECT 21.454 36.795 26.514 36.872 ;
        RECT 21.408 36.841 26.468 36.918 ;
        RECT 21.362 36.887 26.422 36.964 ;
        RECT 21.316 36.933 26.376 37.01 ;
        RECT 21.27 36.979 26.33 37.056 ;
        RECT 21.224 37.025 26.284 37.102 ;
        RECT 21.178 37.071 26.238 37.148 ;
        RECT 21.132 37.117 26.192 37.194 ;
        RECT 21.086 37.163 26.146 37.24 ;
        RECT 21.04 37.209 26.1 37.286 ;
        RECT 20.994 37.255 26.054 37.332 ;
        RECT 20.948 37.301 26.008 37.378 ;
        RECT 20.902 37.347 25.962 37.424 ;
        RECT 20.856 37.393 25.916 37.47 ;
        RECT 20.81 37.439 25.87 37.516 ;
        RECT 20.764 37.485 25.824 37.562 ;
        RECT 20.718 37.531 25.778 37.608 ;
        RECT 20.672 37.577 25.732 37.654 ;
        RECT 20.626 37.623 25.686 37.7 ;
        RECT 20.58 37.669 25.64 37.746 ;
        RECT 20.534 37.715 25.594 37.792 ;
        RECT 20.488 37.761 25.548 37.838 ;
        RECT 20.442 37.807 25.502 37.884 ;
        RECT 20.396 37.853 25.456 37.93 ;
        RECT 20.35 37.899 25.41 37.976 ;
        RECT 20.304 37.945 25.364 38.022 ;
        RECT 20.258 37.991 25.318 38.068 ;
        RECT 20.212 38.037 25.272 38.114 ;
        RECT 20.166 38.083 25.226 38.16 ;
        RECT 20.12 38.129 25.18 38.206 ;
        RECT 20.074 38.175 25.134 38.252 ;
        RECT 20.028 38.221 25.088 38.298 ;
        RECT 19.982 38.267 25.042 38.344 ;
        RECT 19.936 38.313 24.996 38.39 ;
        RECT 19.89 38.359 24.95 38.436 ;
        RECT 19.844 38.405 24.904 38.482 ;
        RECT 19.798 38.451 24.858 38.528 ;
        RECT 19.752 38.497 24.812 38.574 ;
        RECT 19.706 38.543 24.766 38.62 ;
        RECT 19.66 38.589 24.72 38.666 ;
        RECT 19.614 38.635 24.674 38.712 ;
        RECT 19.568 38.681 24.628 38.758 ;
        RECT 19.522 38.727 24.582 38.804 ;
        RECT 19.476 38.773 24.536 38.85 ;
        RECT 19.43 38.819 24.49 38.896 ;
        RECT 19.384 38.865 24.444 38.942 ;
        RECT 19.338 38.911 24.398 38.988 ;
        RECT 19.292 38.957 24.352 39.034 ;
        RECT 19.246 39.003 24.306 39.08 ;
        RECT 19.2 39.049 24.26 39.126 ;
        RECT 19.154 39.095 24.214 39.172 ;
        RECT 19.108 39.141 24.168 39.218 ;
        RECT 19.062 39.187 24.122 39.264 ;
        RECT 19.016 39.233 24.076 39.31 ;
        RECT 18.97 39.279 24.03 39.356 ;
        RECT 18.924 39.325 23.984 39.402 ;
        RECT 18.878 39.371 23.938 39.448 ;
        RECT 18.832 39.417 23.892 39.494 ;
        RECT 18.786 39.463 23.846 39.54 ;
        RECT 18.74 39.509 23.8 39.586 ;
        RECT 18.694 39.555 23.754 39.632 ;
        RECT 18.648 39.601 23.708 39.678 ;
        RECT 18.602 39.647 23.662 39.724 ;
        RECT 18.556 39.693 23.616 39.77 ;
        RECT 18.51 39.739 23.57 39.816 ;
        RECT 18.464 39.785 23.524 39.862 ;
        RECT 18.418 39.831 23.478 39.908 ;
        RECT 18.372 39.877 23.432 39.954 ;
        RECT 18.326 39.923 23.386 40 ;
        RECT 18.28 39.969 23.34 40.046 ;
        RECT 18.234 40.015 23.294 40.092 ;
        RECT 18.188 40.061 23.248 40.138 ;
        RECT 18.142 40.107 23.202 40.184 ;
        RECT 18.096 40.153 23.156 40.23 ;
        RECT 18.05 40.199 23.11 40.276 ;
        RECT 18.004 40.245 23.064 40.322 ;
        RECT 17.958 40.291 23.018 40.368 ;
        RECT 17.912 40.337 22.972 40.414 ;
        RECT 17.866 40.383 22.926 40.46 ;
        RECT 17.82 40.429 22.88 40.506 ;
        RECT 17.774 40.475 22.834 40.552 ;
        RECT 17.728 40.521 22.788 40.598 ;
        RECT 17.682 40.567 22.742 40.644 ;
        RECT 17.636 40.613 22.696 40.69 ;
        RECT 17.59 40.659 22.65 40.736 ;
        RECT 17.544 40.705 22.604 40.782 ;
        RECT 17.498 40.751 22.558 40.828 ;
        RECT 17.452 40.797 22.512 40.874 ;
        RECT 17.406 40.843 22.466 40.92 ;
        RECT 17.36 40.889 22.42 40.966 ;
        RECT 17.314 40.935 22.374 41.012 ;
        RECT 17.268 40.981 22.328 41.058 ;
        RECT 17.222 41.027 22.282 41.104 ;
        RECT 17.176 41.073 22.236 41.15 ;
        RECT 17.13 41.119 22.19 41.196 ;
        RECT 17.084 41.165 22.144 41.242 ;
        RECT 17.038 41.211 22.098 41.288 ;
        RECT 16.992 41.257 22.052 41.334 ;
        RECT 16.946 41.303 22.006 41.38 ;
        RECT 16.9 41.349 21.96 41.426 ;
        RECT 16.854 41.395 21.914 41.472 ;
        RECT 16.808 41.441 21.868 41.518 ;
        RECT 16.762 41.487 21.822 41.564 ;
        RECT 16.716 41.533 21.776 41.61 ;
        RECT 16.67 41.579 21.73 41.656 ;
        RECT 16.624 41.625 21.684 41.702 ;
        RECT 16.578 41.671 21.638 41.748 ;
        RECT 16.532 41.717 21.592 41.794 ;
        RECT 16.486 41.763 21.546 41.84 ;
        RECT 16.44 41.809 21.5 41.886 ;
        RECT 16.394 41.855 21.454 41.932 ;
        RECT 16.348 41.901 21.408 41.978 ;
        RECT 16.302 41.947 21.362 42.024 ;
        RECT 16.256 41.993 21.316 42.07 ;
        RECT 16.21 42.039 21.27 42.116 ;
        RECT 16.164 42.085 21.224 42.162 ;
        RECT 16.118 42.131 21.178 42.208 ;
        RECT 16.072 42.177 21.132 42.254 ;
        RECT 16.026 42.223 21.086 42.3 ;
        RECT 15.98 42.269 21.04 42.346 ;
        RECT 15.934 42.315 20.994 42.392 ;
        RECT 15.888 42.361 20.948 42.438 ;
        RECT 15.842 42.407 20.902 42.484 ;
        RECT 15.796 42.453 20.856 42.53 ;
        RECT 15.75 42.499 20.81 42.576 ;
        RECT 15.704 42.545 20.764 42.622 ;
        RECT 15.658 42.591 20.718 42.668 ;
        RECT 15.612 42.637 20.672 42.714 ;
        RECT 15.566 42.683 20.626 42.76 ;
        RECT 15.52 42.729 20.58 42.806 ;
        RECT 15.474 42.775 20.534 42.852 ;
        RECT 15.428 42.821 20.488 42.898 ;
        RECT 15.382 42.867 20.442 42.944 ;
        RECT 15.336 42.913 20.396 42.99 ;
        RECT 15.29 42.959 20.35 43.036 ;
        RECT 15.244 43.005 20.304 43.082 ;
        RECT 15.198 43.051 20.258 43.128 ;
        RECT 15.152 43.097 20.212 43.174 ;
        RECT 15.106 43.143 20.166 43.22 ;
        RECT 15.06 43.189 20.12 43.266 ;
        RECT 15.014 43.235 20.074 43.312 ;
        RECT 14.968 43.281 20.028 43.358 ;
        RECT 14.922 43.327 19.982 43.404 ;
        RECT 14.876 43.373 19.936 43.45 ;
        RECT 14.83 43.419 19.89 43.496 ;
        RECT 14.784 43.465 19.844 43.542 ;
        RECT 14.738 43.511 19.798 43.588 ;
        RECT 14.692 43.557 19.752 43.634 ;
        RECT 14.646 43.603 19.706 43.68 ;
        RECT 14.6 43.649 19.66 43.726 ;
        RECT 14.554 43.695 19.614 43.772 ;
        RECT 14.508 43.741 19.568 43.818 ;
        RECT 14.462 43.787 19.522 43.864 ;
        RECT 14.416 43.833 19.476 43.91 ;
        RECT 14.37 43.879 19.43 43.956 ;
        RECT 14.324 43.925 19.384 44.002 ;
        RECT 14.278 43.971 19.338 44.048 ;
        RECT 14.232 44.017 19.292 44.094 ;
        RECT 14.186 44.063 19.246 44.14 ;
        RECT 14.14 44.109 19.2 44.186 ;
        RECT 14.094 44.155 19.154 44.232 ;
        RECT 14.048 44.201 19.108 44.278 ;
        RECT 14.002 44.247 19.062 44.324 ;
        RECT 13.956 44.293 19.016 44.37 ;
        RECT 13.91 44.339 18.97 44.416 ;
        RECT 13.864 44.385 18.924 44.462 ;
        RECT 13.818 44.431 18.878 44.508 ;
        RECT 13.772 44.477 18.832 44.554 ;
        RECT 13.726 44.523 18.786 44.6 ;
        RECT 13.68 44.569 18.74 44.646 ;
        RECT 13.634 44.615 18.694 44.692 ;
        RECT 13.588 44.661 18.648 44.738 ;
        RECT 13.542 44.707 18.602 44.784 ;
        RECT 13.496 44.753 18.556 44.83 ;
        RECT 13.45 44.799 18.51 44.876 ;
        RECT 13.404 44.845 18.464 44.922 ;
        RECT 13.358 44.891 18.418 44.968 ;
        RECT 13.312 44.937 18.372 45.014 ;
        RECT 13.266 44.983 18.326 45.06 ;
        RECT 13.22 45.029 18.28 45.106 ;
        RECT 13.174 45.075 18.234 45.152 ;
        RECT 13.128 45.121 18.188 45.198 ;
        RECT 13.082 45.167 18.142 45.244 ;
        RECT 13.036 45.213 18.096 45.29 ;
        RECT 12.99 45.259 18.05 45.336 ;
        RECT 12.944 45.305 18.004 45.382 ;
        RECT 12.898 45.351 17.958 45.428 ;
        RECT 12.852 45.397 17.912 45.474 ;
        RECT 12.806 45.443 17.866 45.52 ;
        RECT 12.76 45.489 17.82 45.566 ;
        RECT 12.714 45.535 17.774 45.612 ;
        RECT 12.668 45.581 17.728 45.658 ;
        RECT 12.622 45.627 17.682 45.704 ;
        RECT 12.576 45.673 17.636 45.75 ;
        RECT 12.53 45.719 17.59 45.796 ;
        RECT 12.484 45.765 17.544 45.842 ;
        RECT 12.438 45.811 17.498 45.888 ;
        RECT 12.392 45.857 17.452 45.934 ;
        RECT 12.346 45.903 17.406 45.98 ;
        RECT 12.3 45.949 17.36 46.026 ;
        RECT 12.254 45.995 17.314 46.072 ;
        RECT 12.208 46.041 17.268 46.118 ;
        RECT 12.162 46.087 17.222 46.164 ;
        RECT 12.116 46.133 17.176 46.21 ;
        RECT 12.07 46.179 17.13 46.256 ;
        RECT 12.024 46.225 17.084 46.302 ;
        RECT 11.978 46.271 17.038 46.348 ;
        RECT 11.932 46.317 16.992 46.394 ;
        RECT 11.886 46.363 16.946 46.44 ;
        RECT 11.84 46.409 16.9 46.486 ;
        RECT 11.794 46.455 16.854 46.532 ;
        RECT 11.748 46.501 16.808 46.578 ;
        RECT 11.702 46.547 16.762 46.624 ;
        RECT 11.656 46.593 16.716 46.67 ;
        RECT 11.61 46.639 16.67 46.716 ;
        RECT 11.564 46.685 16.624 46.762 ;
        RECT 11.518 46.731 16.578 46.808 ;
        RECT 11.472 46.777 16.532 46.854 ;
        RECT 11.426 46.823 16.486 46.9 ;
        RECT 11.38 46.869 16.44 46.946 ;
        RECT 11.334 46.915 16.394 46.992 ;
        RECT 11.288 46.961 16.348 47.038 ;
        RECT 11.242 47.007 16.302 47.084 ;
        RECT 11.196 47.053 16.256 47.13 ;
        RECT 11.15 47.099 16.21 47.176 ;
        RECT 11.104 47.145 16.164 47.222 ;
        RECT 11.058 47.191 16.118 47.268 ;
        RECT 11.012 47.237 16.072 47.314 ;
        RECT 10.966 47.283 16.026 47.36 ;
        RECT 10.92 47.329 15.98 47.406 ;
        RECT 10.874 47.375 15.934 47.452 ;
        RECT 10.828 47.421 15.888 47.498 ;
        RECT 10.782 47.467 15.842 47.544 ;
        RECT 10.736 47.513 15.796 47.59 ;
        RECT 10.69 47.559 15.75 47.636 ;
        RECT 10.644 47.605 15.704 47.682 ;
        RECT 10.598 47.651 15.658 47.728 ;
        RECT 10.552 47.697 15.612 47.774 ;
        RECT 10.506 47.743 15.566 47.82 ;
        RECT 10.46 47.789 15.52 47.866 ;
        RECT 10.414 47.835 15.474 47.912 ;
        RECT 10.368 47.881 15.428 47.958 ;
        RECT 10.322 47.927 15.382 48.004 ;
        RECT 10.276 47.973 15.336 48.05 ;
        RECT 10.23 48.019 15.29 48.096 ;
        RECT 10.184 48.065 15.244 48.142 ;
        RECT 10.138 48.111 15.198 48.188 ;
        RECT 10.092 48.157 15.152 48.234 ;
        RECT 10.046 48.203 15.106 48.28 ;
        RECT 10 48.249 15.06 48.326 ;
        RECT 9.954 48.295 15.014 48.372 ;
        RECT 9.908 48.341 14.968 48.418 ;
        RECT 9.862 48.387 14.922 48.464 ;
        RECT 9.816 48.433 14.876 48.51 ;
        RECT 9.77 48.479 14.83 48.556 ;
        RECT 9.724 48.525 14.784 48.602 ;
        RECT 9.678 48.571 14.738 48.648 ;
        RECT 9.632 48.617 14.692 48.694 ;
        RECT 9.586 48.663 14.646 48.74 ;
        RECT 9.54 48.709 14.6 48.786 ;
        RECT 9.494 48.755 14.554 48.832 ;
        RECT 9.448 48.801 14.508 48.878 ;
        RECT 9.402 48.847 14.462 48.924 ;
        RECT 9.356 48.893 14.416 48.97 ;
        RECT 9.31 48.939 14.37 49.016 ;
        RECT 9.264 48.985 14.324 49.062 ;
        RECT 9.218 49.031 14.278 49.108 ;
        RECT 9.172 49.077 14.232 49.154 ;
        RECT 9.126 49.123 14.186 49.2 ;
        RECT 9.08 49.169 14.14 49.246 ;
        RECT 9.034 49.215 14.094 49.292 ;
        RECT 8.988 49.261 14.048 49.338 ;
        RECT 8.942 49.307 14.002 49.384 ;
        RECT 8.896 49.353 13.956 49.43 ;
        RECT 8.85 49.399 13.91 49.476 ;
        RECT 8.804 49.445 13.864 49.522 ;
        RECT 8.758 49.491 13.818 49.568 ;
        RECT 8.712 49.537 13.772 49.614 ;
    END
    PORT
      LAYER IB ;
        RECT 58.414 26.45 80 30.05 ;
        RECT 54.798 30.043 59.905 30.06 ;
        RECT 53.372 31.469 58.46 31.518 ;
        RECT 58.386 26.464 58.414 31.555 ;
        RECT 53.326 31.515 58.386 31.592 ;
        RECT 53.418 31.423 58.506 31.472 ;
        RECT 58.34 26.501 58.386 31.592 ;
        RECT 53.28 31.561 58.34 31.638 ;
        RECT 53.464 31.377 58.552 31.426 ;
        RECT 58.294 26.547 58.34 31.638 ;
        RECT 53.234 31.607 58.294 31.684 ;
        RECT 53.51 31.331 58.598 31.38 ;
        RECT 58.248 26.593 58.294 31.684 ;
        RECT 53.188 31.653 58.248 31.73 ;
        RECT 53.556 31.285 58.644 31.334 ;
        RECT 58.202 26.639 58.248 31.73 ;
        RECT 53.142 31.699 58.202 31.776 ;
        RECT 53.602 31.239 58.69 31.288 ;
        RECT 58.156 26.685 58.202 31.776 ;
        RECT 53.096 31.745 58.156 31.822 ;
        RECT 53.648 31.193 58.736 31.242 ;
        RECT 58.11 26.731 58.156 31.822 ;
        RECT 53.05 31.791 58.11 31.868 ;
        RECT 53.694 31.147 58.782 31.196 ;
        RECT 58.064 26.777 58.11 31.868 ;
        RECT 53.004 31.837 58.064 31.914 ;
        RECT 53.74 31.101 58.828 31.15 ;
        RECT 58.018 26.823 58.064 31.914 ;
        RECT 52.958 31.883 58.018 31.96 ;
        RECT 53.786 31.055 58.874 31.104 ;
        RECT 57.972 26.869 58.018 31.96 ;
        RECT 52.912 31.929 57.972 32.006 ;
        RECT 53.832 31.009 58.92 31.058 ;
        RECT 57.926 26.915 57.972 32.006 ;
        RECT 52.866 31.975 57.926 32.052 ;
        RECT 53.878 30.963 58.966 31.012 ;
        RECT 57.88 26.961 57.926 32.052 ;
        RECT 52.82 32.021 57.88 32.098 ;
        RECT 53.924 30.917 59.012 30.966 ;
        RECT 57.834 27.007 57.88 32.098 ;
        RECT 52.774 32.067 57.834 32.144 ;
        RECT 53.97 30.871 59.058 30.92 ;
        RECT 57.788 27.053 57.834 32.144 ;
        RECT 52.728 32.113 57.788 32.19 ;
        RECT 54.016 30.825 59.104 30.874 ;
        RECT 57.742 27.099 57.788 32.19 ;
        RECT 52.682 32.159 57.742 32.236 ;
        RECT 54.062 30.779 59.15 30.828 ;
        RECT 57.696 27.145 57.742 32.236 ;
        RECT 52.636 32.205 57.696 32.282 ;
        RECT 54.108 30.733 59.196 30.782 ;
        RECT 57.65 27.191 57.696 32.282 ;
        RECT 52.59 32.251 57.65 32.328 ;
        RECT 54.154 30.687 59.242 30.736 ;
        RECT 57.604 27.237 57.65 32.328 ;
        RECT 52.544 32.297 57.604 32.374 ;
        RECT 54.2 30.641 59.288 30.69 ;
        RECT 57.558 27.283 57.604 32.374 ;
        RECT 52.498 32.343 57.558 32.42 ;
        RECT 54.246 30.595 59.334 30.644 ;
        RECT 57.512 27.329 57.558 32.42 ;
        RECT 52.452 32.389 57.512 32.466 ;
        RECT 54.292 30.549 59.38 30.598 ;
        RECT 57.466 27.375 57.512 32.466 ;
        RECT 52.406 32.435 57.466 32.512 ;
        RECT 54.338 30.503 59.426 30.552 ;
        RECT 57.42 27.421 57.466 32.512 ;
        RECT 52.36 32.481 57.42 32.558 ;
        RECT 54.384 30.457 59.472 30.506 ;
        RECT 57.374 27.467 57.42 32.558 ;
        RECT 52.314 32.527 57.374 32.604 ;
        RECT 54.43 30.411 59.518 30.46 ;
        RECT 57.328 27.513 57.374 32.604 ;
        RECT 52.268 32.573 57.328 32.65 ;
        RECT 54.476 30.365 59.564 30.414 ;
        RECT 57.282 27.559 57.328 32.65 ;
        RECT 52.222 32.619 57.282 32.696 ;
        RECT 54.522 30.319 59.61 30.368 ;
        RECT 57.236 27.605 57.282 32.696 ;
        RECT 52.176 32.665 57.236 32.742 ;
        RECT 54.568 30.273 59.656 30.322 ;
        RECT 57.19 27.651 57.236 32.742 ;
        RECT 52.13 32.711 57.19 32.788 ;
        RECT 54.614 30.227 59.702 30.276 ;
        RECT 57.144 27.697 57.19 32.788 ;
        RECT 52.084 32.757 57.144 32.834 ;
        RECT 54.66 30.181 59.748 30.23 ;
        RECT 57.098 27.743 57.144 32.834 ;
        RECT 52.038 32.803 57.098 32.88 ;
        RECT 54.706 30.135 59.794 30.184 ;
        RECT 57.052 27.789 57.098 32.88 ;
        RECT 51.992 32.849 57.052 32.926 ;
        RECT 54.752 30.089 59.84 30.138 ;
        RECT 57.006 27.835 57.052 32.926 ;
        RECT 51.946 32.895 57.006 32.972 ;
        RECT 54.798 30.043 59.886 30.092 ;
        RECT 56.96 27.881 57.006 32.972 ;
        RECT 51.9 32.941 56.96 33.018 ;
        RECT 54.844 29.997 80 30.05 ;
        RECT 56.914 27.927 56.96 33.018 ;
        RECT 51.854 32.987 56.914 33.064 ;
        RECT 54.89 29.951 80 30.05 ;
        RECT 56.868 27.973 56.914 33.064 ;
        RECT 51.808 33.033 56.868 33.11 ;
        RECT 54.936 29.905 80 30.05 ;
        RECT 56.822 28.019 56.868 33.11 ;
        RECT 51.762 33.079 56.822 33.156 ;
        RECT 54.982 29.859 80 30.05 ;
        RECT 56.776 28.065 56.822 33.156 ;
        RECT 51.716 33.125 56.776 33.202 ;
        RECT 55.028 29.813 80 30.05 ;
        RECT 56.73 28.111 56.776 33.202 ;
        RECT 51.67 33.171 56.73 33.248 ;
        RECT 55.074 29.767 80 30.05 ;
        RECT 56.684 28.157 56.73 33.248 ;
        RECT 51.624 33.217 56.684 33.294 ;
        RECT 55.12 29.721 80 30.05 ;
        RECT 56.638 28.203 56.684 33.294 ;
        RECT 51.578 33.263 56.638 33.34 ;
        RECT 55.166 29.675 80 30.05 ;
        RECT 56.592 28.249 56.638 33.34 ;
        RECT 51.532 33.309 56.592 33.386 ;
        RECT 55.212 29.629 80 30.05 ;
        RECT 56.546 28.295 56.592 33.386 ;
        RECT 51.486 33.355 56.546 33.432 ;
        RECT 55.258 29.583 80 30.05 ;
        RECT 56.5 28.341 56.546 33.432 ;
        RECT 51.44 33.401 56.5 33.478 ;
        RECT 55.304 29.537 80 30.05 ;
        RECT 56.454 28.387 56.5 33.478 ;
        RECT 51.394 33.447 56.454 33.524 ;
        RECT 55.35 29.491 80 30.05 ;
        RECT 56.408 28.433 56.454 33.524 ;
        RECT 51.348 33.493 56.408 33.57 ;
        RECT 55.396 29.445 80 30.05 ;
        RECT 56.362 28.479 56.408 33.57 ;
        RECT 51.302 33.539 56.362 33.616 ;
        RECT 55.442 29.399 80 30.05 ;
        RECT 56.316 28.525 56.362 33.616 ;
        RECT 51.256 33.585 56.316 33.662 ;
        RECT 55.488 29.353 80 30.05 ;
        RECT 56.27 28.571 56.316 33.662 ;
        RECT 51.21 33.631 56.27 33.708 ;
        RECT 55.534 29.307 80 30.05 ;
        RECT 56.224 28.617 56.27 33.708 ;
        RECT 51.164 33.677 56.224 33.754 ;
        RECT 55.58 29.261 80 30.05 ;
        RECT 56.178 28.663 56.224 33.754 ;
        RECT 51.118 33.723 56.178 33.8 ;
        RECT 55.626 29.215 80 30.05 ;
        RECT 56.132 28.709 56.178 33.8 ;
        RECT 51.072 33.769 56.132 33.846 ;
        RECT 55.672 29.169 80 30.05 ;
        RECT 56.086 28.755 56.132 33.846 ;
        RECT 51.026 33.815 56.086 33.892 ;
        RECT 55.718 29.123 80 30.05 ;
        RECT 56.04 28.801 56.086 33.892 ;
        RECT 50.98 33.861 56.04 33.938 ;
        RECT 55.764 29.077 80 30.05 ;
        RECT 55.994 28.847 56.04 33.938 ;
        RECT 50.934 33.907 55.994 33.984 ;
        RECT 55.81 29.031 80 30.05 ;
        RECT 55.948 28.893 55.994 33.984 ;
        RECT 50.888 33.953 55.948 34.03 ;
        RECT 55.856 28.985 80 30.05 ;
        RECT 55.902 28.939 55.948 34.03 ;
        RECT 50.842 33.999 55.902 34.076 ;
        RECT 50.796 34.045 55.856 34.122 ;
        RECT 50.75 34.091 55.81 34.168 ;
        RECT 50.704 34.137 55.764 34.214 ;
        RECT 50.658 34.183 55.718 34.26 ;
        RECT 50.612 34.229 55.672 34.306 ;
        RECT 50.566 34.275 55.626 34.352 ;
        RECT 50.52 34.321 55.58 34.398 ;
        RECT 50.474 34.367 55.534 34.444 ;
        RECT 50.428 34.413 55.488 34.49 ;
        RECT 50.382 34.459 55.442 34.536 ;
        RECT 50.336 34.505 55.396 34.582 ;
        RECT 50.29 34.551 55.35 34.628 ;
        RECT 50.244 34.597 55.304 34.674 ;
        RECT 50.198 34.643 55.258 34.72 ;
        RECT 50.152 34.689 55.212 34.766 ;
        RECT 50.106 34.735 55.166 34.812 ;
        RECT 50.06 34.781 55.12 34.858 ;
        RECT 50.014 34.827 55.074 34.904 ;
        RECT 49.968 34.873 55.028 34.95 ;
        RECT 49.922 34.919 54.982 34.996 ;
        RECT 49.876 34.965 54.936 35.042 ;
        RECT 49.83 35.011 54.89 35.088 ;
        RECT 49.784 35.057 54.844 35.134 ;
        RECT 49.738 35.103 54.798 35.18 ;
        RECT 49.692 35.149 54.752 35.226 ;
        RECT 49.646 35.195 54.706 35.272 ;
        RECT 49.6 35.241 54.66 35.318 ;
        RECT 49.554 35.287 54.614 35.364 ;
        RECT 49.508 35.333 54.568 35.41 ;
        RECT 49.462 35.379 54.522 35.456 ;
        RECT 49.416 35.425 54.476 35.502 ;
        RECT 49.37 35.471 54.43 35.548 ;
        RECT 49.324 35.517 54.384 35.594 ;
        RECT 49.278 35.563 54.338 35.64 ;
        RECT 49.232 35.609 54.292 35.686 ;
        RECT 49.186 35.655 54.246 35.732 ;
        RECT 49.14 35.701 54.2 35.778 ;
        RECT 49.094 35.747 54.154 35.824 ;
        RECT 49.048 35.793 54.108 35.87 ;
        RECT 49.002 35.839 54.062 35.916 ;
        RECT 48.956 35.885 54.016 35.962 ;
        RECT 48.91 35.931 53.97 36.008 ;
        RECT 48.864 35.977 53.924 36.054 ;
        RECT 48.818 36.023 53.878 36.1 ;
        RECT 48.772 36.069 53.832 36.146 ;
        RECT 48.726 36.115 53.786 36.192 ;
        RECT 48.68 36.161 53.74 36.238 ;
        RECT 48.634 36.207 53.694 36.284 ;
        RECT 48.588 36.253 53.648 36.33 ;
        RECT 48.542 36.299 53.602 36.376 ;
        RECT 48.496 36.345 53.556 36.422 ;
        RECT 48.45 36.391 53.51 36.468 ;
        RECT 48.404 36.437 53.464 36.514 ;
        RECT 48.358 36.483 53.418 36.56 ;
        RECT 48.312 36.529 53.372 36.606 ;
        RECT 48.266 36.575 53.326 36.652 ;
        RECT 48.22 36.621 53.28 36.698 ;
        RECT 48.174 36.667 53.234 36.744 ;
        RECT 48.128 36.713 53.188 36.79 ;
        RECT 48.082 36.759 53.142 36.836 ;
        RECT 48.036 36.805 53.096 36.882 ;
        RECT 47.99 36.851 53.05 36.928 ;
        RECT 47.944 36.897 53.004 36.974 ;
        RECT 47.898 36.943 52.958 37.02 ;
        RECT 47.852 36.989 52.912 37.066 ;
        RECT 47.806 37.035 52.866 37.112 ;
        RECT 47.76 37.081 52.82 37.158 ;
        RECT 47.714 37.127 52.774 37.204 ;
        RECT 47.668 37.173 52.728 37.25 ;
        RECT 47.622 37.219 52.682 37.296 ;
        RECT 47.576 37.265 52.636 37.342 ;
        RECT 47.53 37.311 52.59 37.388 ;
        RECT 47.484 37.357 52.544 37.434 ;
        RECT 47.438 37.403 52.498 37.48 ;
        RECT 47.392 37.449 52.452 37.526 ;
        RECT 47.346 37.495 52.406 37.572 ;
        RECT 47.3 37.541 52.36 37.618 ;
        RECT 47.254 37.587 52.314 37.664 ;
        RECT 47.208 37.633 52.268 37.71 ;
        RECT 47.162 37.679 52.222 37.756 ;
        RECT 47.116 37.725 52.176 37.802 ;
        RECT 47.07 37.771 52.13 37.848 ;
        RECT 47.024 37.817 52.084 37.894 ;
        RECT 46.978 37.863 52.038 37.94 ;
        RECT 46.932 37.909 51.992 37.986 ;
        RECT 46.886 37.955 51.946 38.032 ;
        RECT 46.84 38.001 51.9 38.078 ;
        RECT 46.794 38.047 51.854 38.124 ;
        RECT 46.748 38.093 51.808 38.17 ;
        RECT 46.702 38.139 51.762 38.216 ;
        RECT 46.656 38.185 51.716 38.262 ;
        RECT 46.61 38.231 51.67 38.308 ;
        RECT 46.564 38.277 51.624 38.354 ;
        RECT 46.518 38.323 51.578 38.4 ;
        RECT 46.472 38.369 51.532 38.446 ;
        RECT 46.426 38.415 51.486 38.492 ;
        RECT 46.38 38.461 51.44 38.538 ;
        RECT 46.334 38.507 51.394 38.584 ;
        RECT 46.288 38.553 51.348 38.63 ;
        RECT 46.242 38.599 51.302 38.676 ;
        RECT 46.196 38.645 51.256 38.722 ;
        RECT 46.15 38.691 51.21 38.768 ;
        RECT 46.104 38.737 51.164 38.814 ;
        RECT 46.058 38.783 51.118 38.86 ;
        RECT 46.012 38.829 51.072 38.906 ;
        RECT 45.966 38.875 51.026 38.952 ;
        RECT 45.92 38.921 50.98 38.998 ;
        RECT 45.874 38.967 50.934 39.044 ;
        RECT 45.828 39.013 50.888 39.09 ;
        RECT 45.782 39.059 50.842 39.136 ;
        RECT 45.736 39.105 50.796 39.182 ;
        RECT 45.69 39.151 50.75 39.228 ;
        RECT 45.644 39.197 50.704 39.274 ;
        RECT 45.598 39.243 50.658 39.32 ;
        RECT 45.552 39.289 50.612 39.366 ;
        RECT 45.506 39.335 50.566 39.412 ;
        RECT 45.46 39.381 50.52 39.458 ;
        RECT 45.414 39.427 50.474 39.504 ;
        RECT 45.368 39.473 50.428 39.55 ;
        RECT 45.322 39.519 50.382 39.596 ;
        RECT 45.276 39.565 50.336 39.642 ;
        RECT 45.23 39.611 50.29 39.688 ;
        RECT 45.184 39.657 50.244 39.734 ;
        RECT 45.138 39.703 50.198 39.78 ;
        RECT 45.092 39.749 50.152 39.826 ;
        RECT 45.046 39.795 50.106 39.872 ;
        RECT 45 39.841 50.06 39.918 ;
        RECT 44.954 39.887 50.014 39.964 ;
        RECT 44.908 39.933 49.968 40.01 ;
        RECT 44.862 39.979 49.922 40.056 ;
        RECT 44.816 40.025 49.876 40.102 ;
        RECT 44.77 40.071 49.83 40.148 ;
        RECT 44.724 40.117 49.784 40.194 ;
        RECT 44.678 40.163 49.738 40.24 ;
        RECT 44.632 40.209 49.692 40.286 ;
        RECT 44.586 40.255 49.646 40.332 ;
        RECT 44.54 40.301 49.6 40.378 ;
        RECT 44.494 40.347 49.554 40.424 ;
        RECT 44.448 40.393 49.508 40.47 ;
        RECT 44.402 40.439 49.462 40.516 ;
        RECT 44.356 40.485 49.416 40.562 ;
        RECT 44.31 40.531 49.37 40.608 ;
        RECT 44.264 40.577 49.324 40.654 ;
        RECT 44.218 40.623 49.278 40.7 ;
        RECT 44.172 40.669 49.232 40.746 ;
        RECT 44.126 40.715 49.186 40.792 ;
        RECT 44.08 40.761 49.14 40.838 ;
        RECT 44.034 40.807 49.094 40.884 ;
        RECT 43.988 40.853 49.048 40.93 ;
        RECT 43.942 40.899 49.002 40.976 ;
        RECT 43.896 40.945 48.956 41.022 ;
        RECT 43.85 40.991 48.91 41.068 ;
        RECT 43.804 41.037 48.864 41.114 ;
        RECT 43.758 41.083 48.818 41.16 ;
        RECT 43.712 41.129 48.772 41.206 ;
        RECT 43.666 41.175 48.726 41.252 ;
        RECT 43.62 41.221 48.68 41.298 ;
        RECT 43.574 41.267 48.634 41.344 ;
        RECT 43.528 41.313 48.588 41.39 ;
        RECT 43.482 41.359 48.542 41.436 ;
        RECT 43.436 41.405 48.496 41.482 ;
        RECT 43.39 41.451 48.45 41.528 ;
        RECT 43.344 41.497 48.404 41.574 ;
        RECT 43.298 41.543 48.358 41.62 ;
        RECT 43.252 41.589 48.312 41.666 ;
        RECT 43.206 41.635 48.266 41.712 ;
        RECT 43.16 41.681 48.22 41.758 ;
        RECT 43.114 41.727 48.174 41.804 ;
        RECT 43.068 41.773 48.128 41.85 ;
        RECT 43.022 41.819 48.082 41.896 ;
        RECT 42.976 41.865 48.036 41.942 ;
        RECT 42.93 41.911 47.99 41.988 ;
        RECT 42.884 41.957 47.944 42.034 ;
        RECT 42.838 42.003 47.898 42.08 ;
        RECT 42.792 42.049 47.852 42.126 ;
        RECT 42.746 42.095 47.806 42.172 ;
        RECT 42.7 42.141 47.76 42.218 ;
        RECT 42.654 42.187 47.714 42.264 ;
        RECT 42.608 42.233 47.668 42.31 ;
        RECT 42.562 42.279 47.622 42.356 ;
        RECT 42.516 42.325 47.576 42.402 ;
        RECT 42.47 42.371 47.53 42.448 ;
        RECT 42.424 42.417 47.484 42.494 ;
        RECT 42.378 42.463 47.438 42.54 ;
        RECT 42.332 42.509 47.392 42.586 ;
        RECT 42.286 42.555 47.346 42.632 ;
        RECT 42.24 42.601 47.3 42.678 ;
        RECT 42.194 42.647 47.254 42.724 ;
        RECT 42.148 42.693 47.208 42.77 ;
        RECT 42.102 42.739 47.162 42.816 ;
        RECT 42.056 42.785 47.116 42.862 ;
        RECT 42.01 42.831 47.07 42.908 ;
        RECT 41.964 42.877 47.024 42.954 ;
        RECT 41.918 42.923 46.978 43 ;
        RECT 41.872 42.969 46.932 43.046 ;
        RECT 41.826 43.015 46.886 43.092 ;
        RECT 41.78 43.061 46.84 43.138 ;
        RECT 41.734 43.107 46.794 43.184 ;
        RECT 41.688 43.153 46.748 43.23 ;
        RECT 41.642 43.199 46.702 43.276 ;
        RECT 41.596 43.245 46.656 43.322 ;
        RECT 41.55 43.291 46.61 43.368 ;
        RECT 41.504 43.337 46.564 43.414 ;
        RECT 41.458 43.383 46.518 43.46 ;
        RECT 41.412 43.429 46.472 43.506 ;
        RECT 41.366 43.475 46.426 43.552 ;
        RECT 41.32 43.521 46.38 43.598 ;
        RECT 41.274 43.567 46.334 43.644 ;
        RECT 41.228 43.613 46.288 43.69 ;
        RECT 41.182 43.659 46.242 43.736 ;
        RECT 41.136 43.705 46.196 43.782 ;
        RECT 41.09 43.751 46.15 43.828 ;
        RECT 41.044 43.797 46.104 43.874 ;
        RECT 40.998 43.843 46.058 43.92 ;
        RECT 40.952 43.889 46.012 43.966 ;
        RECT 40.906 43.935 45.966 44.012 ;
        RECT 40.86 43.981 45.92 44.058 ;
        RECT 40.814 44.027 45.874 44.104 ;
        RECT 40.768 44.073 45.828 44.15 ;
        RECT 40.722 44.119 45.782 44.196 ;
        RECT 40.676 44.165 45.736 44.242 ;
        RECT 40.63 44.211 45.69 44.288 ;
        RECT 40.584 44.257 45.644 44.334 ;
        RECT 40.538 44.303 45.598 44.38 ;
        RECT 40.492 44.349 45.552 44.426 ;
        RECT 40.446 44.395 45.506 44.472 ;
        RECT 40.4 44.441 45.46 44.518 ;
        RECT 40.354 44.487 45.414 44.564 ;
        RECT 40.308 44.533 45.368 44.61 ;
        RECT 40.262 44.579 45.322 44.656 ;
        RECT 40.216 44.625 45.276 44.702 ;
        RECT 40.17 44.671 45.23 44.748 ;
        RECT 40.124 44.717 45.184 44.794 ;
        RECT 40.078 44.763 45.138 44.84 ;
        RECT 40.032 44.809 45.092 44.886 ;
        RECT 39.986 44.855 45.046 44.932 ;
        RECT 39.94 44.901 45 44.978 ;
        RECT 39.894 44.947 44.954 45.024 ;
        RECT 39.848 44.993 44.908 45.07 ;
        RECT 39.802 45.039 44.862 45.116 ;
        RECT 39.756 45.085 44.816 45.162 ;
        RECT 39.71 45.131 44.77 45.208 ;
        RECT 39.664 45.177 44.724 45.254 ;
        RECT 39.618 45.223 44.678 45.3 ;
        RECT 39.572 45.269 44.632 45.346 ;
        RECT 39.526 45.315 44.586 45.392 ;
        RECT 39.48 45.361 44.54 45.438 ;
        RECT 39.434 45.407 44.494 45.484 ;
        RECT 39.388 45.453 44.448 45.53 ;
        RECT 39.342 45.499 44.402 45.576 ;
        RECT 39.296 45.545 44.356 45.622 ;
        RECT 39.25 45.591 44.31 45.668 ;
        RECT 39.204 45.637 44.264 45.714 ;
        RECT 39.158 45.683 44.218 45.76 ;
        RECT 39.112 45.729 44.172 45.806 ;
        RECT 39.066 45.775 44.126 45.852 ;
        RECT 39.02 45.821 44.08 45.898 ;
        RECT 38.974 45.867 44.034 45.944 ;
        RECT 38.928 45.913 43.988 45.99 ;
        RECT 38.882 45.959 43.942 46.036 ;
        RECT 38.836 46.005 43.896 46.082 ;
        RECT 38.79 46.051 43.85 46.128 ;
        RECT 38.744 46.097 43.804 46.174 ;
        RECT 38.698 46.143 43.758 46.22 ;
        RECT 38.652 46.189 43.712 46.266 ;
        RECT 38.606 46.235 43.666 46.312 ;
        RECT 38.56 46.281 43.62 46.358 ;
        RECT 38.514 46.327 43.574 46.404 ;
        RECT 38.468 46.373 43.528 46.45 ;
        RECT 38.422 46.419 43.482 46.496 ;
        RECT 38.376 46.465 43.436 46.542 ;
        RECT 38.33 46.511 43.39 46.588 ;
        RECT 38.284 46.557 43.344 46.634 ;
        RECT 38.238 46.603 43.298 46.68 ;
        RECT 38.192 46.649 43.252 46.726 ;
        RECT 38.146 46.695 43.206 46.772 ;
        RECT 38.1 46.741 43.16 46.818 ;
        RECT 38.054 46.787 43.114 46.864 ;
        RECT 38.008 46.833 43.068 46.91 ;
        RECT 37.962 46.879 43.022 46.956 ;
        RECT 37.916 46.925 42.976 47.002 ;
        RECT 37.87 46.971 42.93 47.048 ;
        RECT 37.824 47.017 42.884 47.094 ;
        RECT 37.778 47.063 42.838 47.14 ;
        RECT 37.732 47.109 42.792 47.186 ;
        RECT 37.686 47.155 42.746 47.232 ;
        RECT 37.64 47.201 42.7 47.278 ;
        RECT 37.594 47.247 42.654 47.324 ;
        RECT 37.548 47.293 42.608 47.37 ;
        RECT 37.502 47.339 42.562 47.416 ;
        RECT 37.456 47.385 42.516 47.462 ;
        RECT 37.41 47.431 42.47 47.508 ;
        RECT 37.364 47.477 42.424 47.554 ;
        RECT 37.318 47.523 42.378 47.6 ;
        RECT 37.272 47.569 42.332 47.646 ;
        RECT 37.226 47.615 42.286 47.692 ;
        RECT 37.18 47.661 42.24 47.738 ;
        RECT 37.134 47.707 42.194 47.784 ;
        RECT 37.088 47.753 42.148 47.83 ;
        RECT 37.042 47.799 42.102 47.876 ;
        RECT 36.996 47.845 42.056 47.922 ;
        RECT 36.95 47.891 42.01 47.968 ;
        RECT 36.904 47.937 41.964 48.014 ;
        RECT 36.858 47.983 41.918 48.06 ;
        RECT 36.812 48.029 41.872 48.106 ;
        RECT 36.766 48.075 41.826 48.152 ;
        RECT 36.72 48.121 41.78 48.198 ;
        RECT 36.674 48.167 41.734 48.244 ;
        RECT 36.628 48.213 41.688 48.29 ;
        RECT 36.582 48.259 41.642 48.336 ;
        RECT 36.536 48.305 41.596 48.382 ;
        RECT 36.49 48.351 41.55 48.428 ;
        RECT 36.444 48.397 41.504 48.474 ;
        RECT 36.398 48.443 41.458 48.52 ;
        RECT 36.352 48.489 41.412 48.566 ;
        RECT 36.306 48.535 41.366 48.612 ;
        RECT 36.26 48.581 41.32 48.658 ;
        RECT 36.214 48.627 41.274 48.704 ;
        RECT 36.168 48.673 41.228 48.75 ;
        RECT 36.122 48.719 41.182 48.796 ;
        RECT 36.076 48.765 41.136 48.842 ;
        RECT 36.03 48.811 41.09 48.888 ;
        RECT 35.984 48.857 41.044 48.934 ;
        RECT 35.938 48.903 40.998 48.98 ;
        RECT 35.892 48.949 40.952 49.026 ;
        RECT 35.846 48.995 40.906 49.072 ;
        RECT 35.8 49.041 40.86 49.118 ;
        RECT 35.754 49.087 40.814 49.164 ;
        RECT 35.708 49.133 40.768 49.21 ;
        RECT 35.662 49.179 40.722 49.256 ;
        RECT 35.616 49.225 40.676 49.302 ;
        RECT 35.57 49.271 40.63 49.348 ;
        RECT 35.524 49.317 40.584 49.394 ;
        RECT 35.478 49.363 40.538 49.44 ;
        RECT 35.432 49.409 40.492 49.486 ;
        RECT 35.386 49.455 40.446 49.532 ;
        RECT 35.34 49.501 40.4 49.578 ;
        RECT 35.294 49.547 40.354 49.624 ;
        RECT 35.248 49.593 40.308 49.67 ;
        RECT 35.202 49.639 40.262 49.716 ;
        RECT 35.156 49.685 40.216 49.762 ;
        RECT 35.11 49.731 40.17 49.808 ;
        RECT 35.064 49.777 40.124 49.854 ;
        RECT 35.018 49.823 40.078 49.9 ;
        RECT 34.972 49.869 40.032 49.946 ;
        RECT 34.926 49.915 39.986 49.992 ;
        RECT 34.88 49.961 39.94 50.038 ;
        RECT 34.834 50.007 39.894 50.084 ;
        RECT 34.788 50.053 39.848 50.13 ;
        RECT 34.742 50.099 39.802 50.176 ;
        RECT 34.696 50.145 39.756 50.222 ;
        RECT 34.65 50.191 39.71 50.268 ;
        RECT 34.604 50.237 39.664 50.314 ;
        RECT 34.558 50.283 39.618 50.36 ;
        RECT 34.512 50.329 39.572 50.406 ;
        RECT 34.466 50.375 39.526 50.452 ;
        RECT 34.42 50.421 39.48 50.498 ;
        RECT 34.374 50.467 39.434 50.544 ;
        RECT 34.328 50.513 39.388 50.59 ;
        RECT 34.282 50.559 39.342 50.636 ;
        RECT 34.236 50.605 39.296 50.682 ;
        RECT 34.19 50.651 39.25 50.728 ;
        RECT 34.144 50.697 39.204 50.774 ;
        RECT 34.098 50.743 39.158 50.82 ;
        RECT 34.052 50.789 39.112 50.866 ;
        RECT 34.006 50.835 39.066 50.912 ;
        RECT 33.96 50.881 39.02 50.958 ;
        RECT 33.914 50.927 38.974 51.004 ;
        RECT 33.868 50.973 38.928 51.05 ;
        RECT 33.822 51.019 38.882 51.096 ;
        RECT 33.776 51.065 38.836 51.142 ;
        RECT 33.73 51.111 38.79 51.188 ;
        RECT 33.684 51.157 38.744 51.234 ;
        RECT 33.638 51.203 38.698 51.28 ;
        RECT 33.592 51.249 38.652 51.326 ;
        RECT 33.546 51.295 38.606 51.372 ;
        RECT 33.5 51.341 38.56 51.418 ;
        RECT 33.454 51.387 38.514 51.464 ;
        RECT 33.408 51.433 38.468 51.51 ;
        RECT 33.362 51.479 38.422 51.556 ;
        RECT 33.316 51.525 38.376 51.602 ;
        RECT 33.27 51.571 38.33 51.648 ;
        RECT 33.224 51.617 38.284 51.694 ;
        RECT 33.178 51.663 38.238 51.74 ;
        RECT 33.132 51.709 38.192 51.786 ;
        RECT 33.086 51.755 38.146 51.832 ;
        RECT 33.04 51.801 38.1 51.878 ;
        RECT 32.994 51.847 38.054 51.924 ;
        RECT 32.948 51.893 38.008 51.97 ;
        RECT 32.902 51.939 37.962 52.016 ;
        RECT 32.856 51.985 37.916 52.062 ;
        RECT 32.81 52.031 37.87 52.108 ;
        RECT 32.764 52.077 37.824 52.154 ;
        RECT 32.718 52.123 37.778 52.2 ;
        RECT 32.672 52.169 37.732 52.246 ;
        RECT 32.626 52.215 37.686 52.292 ;
        RECT 32.58 52.261 37.64 52.338 ;
        RECT 32.534 52.307 37.594 52.384 ;
        RECT 32.488 52.353 37.548 52.43 ;
        RECT 32.442 52.399 37.502 52.476 ;
        RECT 32.396 52.445 37.456 52.522 ;
        RECT 32.35 52.491 37.41 52.568 ;
        RECT 32.304 52.537 37.364 52.614 ;
        RECT 32.258 52.583 37.318 52.66 ;
        RECT 32.212 52.629 37.272 52.706 ;
        RECT 32.166 52.675 37.226 52.752 ;
        RECT 32.12 52.721 37.18 52.798 ;
        RECT 32.074 52.767 37.134 52.844 ;
        RECT 32.028 52.813 37.088 52.89 ;
        RECT 31.982 52.859 37.042 52.936 ;
        RECT 31.936 52.905 36.996 52.982 ;
        RECT 31.89 52.951 36.95 53.028 ;
        RECT 31.844 52.997 36.904 53.074 ;
        RECT 31.798 53.043 36.858 53.12 ;
        RECT 31.752 53.089 36.812 53.166 ;
        RECT 31.706 53.135 36.766 53.212 ;
        RECT 31.66 53.181 36.72 53.258 ;
        RECT 31.614 53.227 36.674 53.304 ;
        RECT 31.568 53.273 36.628 53.35 ;
        RECT 31.522 53.319 36.582 53.396 ;
        RECT 31.476 53.365 36.536 53.442 ;
        RECT 31.43 53.411 36.49 53.488 ;
        RECT 31.384 53.457 36.444 53.534 ;
        RECT 31.338 53.503 36.398 53.58 ;
        RECT 31.292 53.549 36.352 53.626 ;
        RECT 31.246 53.595 36.306 53.672 ;
        RECT 31.2 53.641 36.26 53.718 ;
        RECT 31.154 53.687 36.214 53.764 ;
        RECT 31.108 53.733 36.168 53.81 ;
        RECT 31.062 53.779 36.122 53.856 ;
        RECT 31.016 53.825 36.076 53.902 ;
        RECT 30.97 53.871 36.03 53.948 ;
        RECT 30.924 53.917 35.984 53.994 ;
        RECT 30.878 53.963 35.938 54.04 ;
        RECT 30.832 54.009 35.892 54.086 ;
        RECT 30.786 54.055 35.846 54.132 ;
        RECT 30.74 54.101 35.8 54.178 ;
        RECT 30.694 54.147 35.754 54.224 ;
        RECT 30.648 54.193 35.708 54.27 ;
        RECT 30.602 54.239 35.662 54.316 ;
        RECT 30.556 54.285 35.616 54.362 ;
        RECT 30.51 54.331 35.57 54.408 ;
        RECT 30.464 54.377 35.524 54.454 ;
        RECT 30.418 54.423 35.478 54.5 ;
        RECT 30.372 54.469 35.432 54.546 ;
        RECT 30.326 54.515 35.386 54.592 ;
        RECT 30.28 54.561 35.34 54.638 ;
        RECT 30.234 54.607 35.294 54.684 ;
        RECT 30.188 54.653 35.248 54.73 ;
        RECT 30.142 54.699 35.202 54.776 ;
        RECT 30.05 54.791 35.156 54.822 ;
        RECT 30.096 54.745 35.156 54.822 ;
        RECT 30.038 54.82 35.11 54.868 ;
        RECT 29.992 54.849 35.064 54.914 ;
        RECT 29.946 54.895 35.018 54.96 ;
        RECT 29.9 54.941 34.972 55.006 ;
        RECT 29.854 54.987 34.926 55.052 ;
        RECT 29.808 55.033 34.88 55.098 ;
        RECT 29.762 55.079 34.834 55.144 ;
        RECT 29.716 55.125 34.788 55.19 ;
        RECT 29.67 55.171 34.742 55.236 ;
        RECT 29.624 55.217 34.696 55.282 ;
        RECT 29.578 55.263 34.65 55.328 ;
        RECT 29.532 55.309 34.604 55.374 ;
        RECT 29.486 55.355 34.558 55.42 ;
        RECT 29.44 55.401 34.512 55.466 ;
        RECT 29.394 55.447 34.466 55.512 ;
        RECT 29.348 55.493 34.42 55.558 ;
        RECT 29.302 55.539 34.374 55.604 ;
        RECT 29.256 55.585 34.328 55.65 ;
        RECT 29.21 55.631 34.282 55.696 ;
        RECT 29.164 55.677 34.236 55.742 ;
        RECT 29.118 55.723 34.19 55.788 ;
        RECT 29.072 55.769 34.144 55.834 ;
        RECT 29.026 55.815 34.098 55.88 ;
        RECT 28.98 55.861 34.052 55.926 ;
        RECT 28.934 55.907 34.006 55.972 ;
        RECT 28.888 55.953 33.96 56.018 ;
        RECT 28.842 55.999 33.914 56.064 ;
        RECT 28.796 56.045 33.868 56.11 ;
        RECT 28.75 56.091 33.822 56.156 ;
        RECT 28.704 56.137 33.776 56.202 ;
        RECT 28.658 56.183 33.73 56.248 ;
        RECT 28.612 56.229 33.684 56.294 ;
        RECT 28.566 56.275 33.638 56.34 ;
        RECT 28.52 56.321 33.592 56.386 ;
        RECT 28.474 56.367 33.546 56.432 ;
        RECT 28.428 56.413 33.5 56.478 ;
        RECT 28.382 56.459 33.454 56.524 ;
        RECT 28.336 56.505 33.408 56.57 ;
        RECT 28.29 56.551 33.362 56.616 ;
        RECT 28.244 56.597 33.316 56.662 ;
        RECT 28.198 56.643 33.27 56.708 ;
        RECT 28.152 56.689 33.224 56.754 ;
        RECT 28.106 56.735 33.178 56.8 ;
        RECT 28.06 56.781 33.132 56.846 ;
        RECT 28.014 56.827 33.086 56.892 ;
        RECT 27.968 56.873 33.04 56.938 ;
        RECT 27.922 56.919 32.994 56.984 ;
        RECT 27.876 56.965 32.948 57.03 ;
        RECT 27.83 57.011 32.902 57.076 ;
        RECT 27.784 57.057 32.856 57.122 ;
        RECT 27.738 57.103 32.81 57.168 ;
        RECT 27.692 57.149 32.764 57.214 ;
        RECT 27.646 57.195 32.718 57.26 ;
        RECT 27.6 57.241 32.672 57.306 ;
        RECT 27.554 57.287 32.626 57.352 ;
        RECT 27.508 57.333 32.58 57.398 ;
        RECT 27.462 57.379 32.534 57.444 ;
        RECT 27.416 57.425 32.488 57.49 ;
        RECT 27.37 57.471 32.442 57.536 ;
        RECT 27.324 57.517 32.396 57.582 ;
        RECT 27.278 57.563 32.35 57.628 ;
        RECT 27.232 57.609 32.304 57.674 ;
        RECT 27.186 57.655 32.258 57.72 ;
        RECT 27.14 57.701 32.212 57.766 ;
        RECT 27.094 57.747 32.166 57.812 ;
        RECT 27.048 57.793 32.12 57.858 ;
        RECT 27.002 57.839 32.074 57.904 ;
        RECT 26.956 57.885 32.028 57.95 ;
        RECT 26.91 57.931 31.982 57.996 ;
        RECT 26.864 57.977 31.936 58.042 ;
        RECT 26.818 58.023 31.89 58.088 ;
        RECT 26.772 58.069 31.844 58.134 ;
        RECT 26.726 58.115 31.798 58.18 ;
        RECT 26.68 58.161 31.752 58.226 ;
        RECT 26.634 58.207 31.706 58.272 ;
        RECT 26.588 58.253 31.66 58.318 ;
        RECT 26.542 58.299 31.614 58.364 ;
        RECT 26.496 58.345 31.568 58.41 ;
        RECT 26.45 58.391 31.522 58.456 ;
        RECT 26.45 58.391 31.476 58.502 ;
        RECT 26.45 58.391 31.43 58.548 ;
        RECT 26.45 58.391 31.384 58.594 ;
        RECT 26.45 58.391 31.338 58.64 ;
        RECT 26.45 58.391 31.292 58.686 ;
        RECT 26.45 58.391 31.246 58.732 ;
        RECT 26.45 58.391 31.2 58.778 ;
        RECT 26.45 58.391 31.154 58.824 ;
        RECT 26.45 58.391 31.108 58.87 ;
        RECT 26.45 58.391 31.062 58.916 ;
        RECT 26.45 58.391 31.016 58.962 ;
        RECT 26.45 58.391 30.97 59.008 ;
        RECT 26.45 58.391 30.924 59.054 ;
        RECT 26.45 58.391 30.878 59.1 ;
        RECT 26.45 58.391 30.832 59.146 ;
        RECT 26.45 58.391 30.786 59.192 ;
        RECT 26.45 58.391 30.74 59.238 ;
        RECT 26.45 58.391 30.694 59.284 ;
        RECT 26.45 58.391 30.648 59.33 ;
        RECT 26.45 58.391 30.602 59.376 ;
        RECT 26.45 58.391 30.556 59.422 ;
        RECT 26.45 58.391 30.51 59.468 ;
        RECT 26.45 58.391 30.464 59.514 ;
        RECT 26.45 58.391 30.418 59.56 ;
        RECT 26.45 58.391 30.372 59.606 ;
        RECT 26.45 58.391 30.326 59.652 ;
        RECT 26.45 58.391 30.28 59.698 ;
        RECT 26.45 58.391 30.234 59.744 ;
        RECT 26.45 58.391 30.188 59.79 ;
        RECT 26.45 58.391 30.142 59.836 ;
        RECT 26.45 58.391 30.096 59.882 ;
        RECT 26.45 58.391 30.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 22.536 55.657 27.596 55.734 ;
        RECT 22.49 55.703 27.55 55.78 ;
        RECT 22.444 55.749 27.504 55.826 ;
        RECT 22.398 55.795 27.458 55.872 ;
        RECT 22.352 55.841 27.412 55.918 ;
        RECT 22.306 55.887 27.366 55.964 ;
        RECT 22.26 55.933 27.32 56.01 ;
        RECT 22.214 55.979 27.274 56.056 ;
        RECT 22.168 56.025 27.228 56.102 ;
        RECT 22.122 56.071 27.182 56.148 ;
        RECT 22.076 56.117 27.136 56.194 ;
        RECT 22.03 56.163 27.09 56.24 ;
        RECT 21.984 56.209 27.044 56.286 ;
        RECT 21.938 56.255 26.998 56.332 ;
        RECT 21.892 56.301 26.952 56.378 ;
        RECT 21.846 56.347 26.906 56.424 ;
        RECT 21.8 56.393 26.86 56.47 ;
        RECT 21.754 56.439 26.814 56.516 ;
        RECT 21.708 56.485 26.768 56.562 ;
        RECT 21.662 56.531 26.722 56.608 ;
        RECT 21.616 56.577 26.676 56.654 ;
        RECT 21.57 56.623 26.63 56.7 ;
        RECT 21.524 56.669 26.584 56.746 ;
        RECT 21.478 56.715 26.538 56.792 ;
        RECT 21.432 56.761 26.492 56.838 ;
        RECT 21.386 56.807 26.446 56.884 ;
        RECT 21.34 56.853 26.4 56.93 ;
        RECT 21.294 56.899 26.354 56.976 ;
        RECT 21.248 56.945 26.308 57.022 ;
        RECT 21.202 56.991 26.262 57.068 ;
        RECT 21.156 57.037 26.216 57.114 ;
        RECT 21.11 57.083 26.17 57.16 ;
        RECT 21.064 57.129 26.124 57.206 ;
        RECT 21.018 57.175 26.078 57.252 ;
        RECT 20.972 57.221 26.032 57.298 ;
        RECT 20.926 57.267 25.986 57.344 ;
        RECT 20.88 57.313 25.94 57.39 ;
        RECT 20.834 57.359 25.894 57.436 ;
        RECT 20.788 57.405 25.848 57.482 ;
        RECT 20.742 57.451 25.802 57.528 ;
        RECT 20.65 57.543 25.756 57.574 ;
        RECT 20.696 57.497 25.756 57.574 ;
        RECT 20.638 57.572 25.71 57.62 ;
        RECT 20.592 57.601 25.664 57.666 ;
        RECT 20.546 57.647 25.618 57.712 ;
        RECT 20.5 57.693 25.572 57.758 ;
        RECT 20.454 57.739 25.526 57.804 ;
        RECT 20.408 57.785 25.48 57.85 ;
        RECT 20.362 57.831 25.434 57.896 ;
        RECT 20.316 57.877 25.388 57.942 ;
        RECT 20.27 57.923 25.342 57.988 ;
        RECT 20.224 57.969 25.296 58.034 ;
        RECT 20.178 58.015 25.25 58.08 ;
        RECT 20.132 58.061 25.204 58.126 ;
        RECT 20.086 58.107 25.158 58.172 ;
        RECT 20.04 58.153 25.112 58.218 ;
        RECT 19.994 58.199 25.066 58.264 ;
        RECT 19.948 58.245 25.02 58.31 ;
        RECT 19.902 58.291 24.974 58.356 ;
        RECT 19.856 58.337 24.928 58.402 ;
        RECT 19.81 58.383 24.882 58.448 ;
        RECT 19.764 58.429 24.836 58.494 ;
        RECT 19.718 58.475 24.79 58.54 ;
        RECT 19.672 58.521 24.744 58.586 ;
        RECT 19.626 58.567 24.698 58.632 ;
        RECT 19.58 58.613 24.652 58.678 ;
        RECT 19.534 58.659 24.606 58.724 ;
        RECT 19.488 58.705 24.56 58.77 ;
        RECT 19.442 58.751 24.514 58.816 ;
        RECT 19.396 58.797 24.468 58.862 ;
        RECT 19.35 58.843 24.422 58.908 ;
        RECT 19.304 58.889 24.376 58.954 ;
        RECT 19.258 58.935 24.33 59 ;
        RECT 19.212 58.981 24.284 59.046 ;
        RECT 19.166 59.027 24.238 59.092 ;
        RECT 19.12 59.073 24.192 59.138 ;
        RECT 19.074 59.119 24.146 59.184 ;
        RECT 19.028 59.165 24.1 59.23 ;
        RECT 18.982 59.211 24.054 59.276 ;
        RECT 18.936 59.257 24.008 59.322 ;
        RECT 18.89 59.303 23.962 59.368 ;
        RECT 18.844 59.349 23.916 59.414 ;
        RECT 18.798 59.395 23.87 59.46 ;
        RECT 18.752 59.441 23.824 59.506 ;
        RECT 18.706 59.487 23.778 59.552 ;
        RECT 18.66 59.533 23.732 59.598 ;
        RECT 18.614 59.579 23.686 59.644 ;
        RECT 18.568 59.625 23.64 59.69 ;
        RECT 18.522 59.671 23.594 59.736 ;
        RECT 18.476 59.717 23.548 59.782 ;
        RECT 18.43 59.763 23.502 59.828 ;
        RECT 18.384 59.809 23.456 59.874 ;
        RECT 18.338 59.855 23.41 59.92 ;
        RECT 18.292 59.901 23.364 59.966 ;
        RECT 18.246 59.947 23.318 60.012 ;
        RECT 18.2 59.993 23.272 60.058 ;
        RECT 18.154 60.039 23.226 60.104 ;
        RECT 18.108 60.085 23.18 60.15 ;
        RECT 18.062 60.131 23.134 60.196 ;
        RECT 18.016 60.177 23.088 60.242 ;
        RECT 17.97 60.223 23.042 60.288 ;
        RECT 17.924 60.269 22.996 60.334 ;
        RECT 17.878 60.315 22.95 60.38 ;
        RECT 17.832 60.361 22.904 60.426 ;
        RECT 17.786 60.407 22.858 60.472 ;
        RECT 17.74 60.453 22.812 60.518 ;
        RECT 17.694 60.499 22.766 60.564 ;
        RECT 17.648 60.545 22.72 60.61 ;
        RECT 17.602 60.591 22.674 60.656 ;
        RECT 17.556 60.637 22.628 60.702 ;
        RECT 17.51 60.683 22.582 60.748 ;
        RECT 17.464 60.729 22.536 60.794 ;
        RECT 17.418 60.775 22.49 60.84 ;
        RECT 17.372 60.821 22.444 60.886 ;
        RECT 17.326 60.867 22.398 60.932 ;
        RECT 17.28 60.913 22.352 60.978 ;
        RECT 17.234 60.959 22.306 61.024 ;
        RECT 17.188 61.005 22.26 61.07 ;
        RECT 17.142 61.051 22.214 61.116 ;
        RECT 17.096 61.097 22.168 61.162 ;
        RECT 17.05 61.143 22.122 61.208 ;
        RECT 17.05 61.143 22.076 61.254 ;
        RECT 17.05 61.143 22.03 61.3 ;
        RECT 17.05 61.143 21.984 61.346 ;
        RECT 17.05 61.143 21.938 61.392 ;
        RECT 17.05 61.143 21.892 61.438 ;
        RECT 17.05 61.143 21.846 61.484 ;
        RECT 17.05 61.143 21.8 61.53 ;
        RECT 17.05 61.143 21.754 61.576 ;
        RECT 17.05 61.143 21.708 61.622 ;
        RECT 17.05 61.143 21.662 61.668 ;
        RECT 17.05 61.143 21.616 61.714 ;
        RECT 17.05 61.143 21.57 61.76 ;
        RECT 17.05 61.143 21.524 61.806 ;
        RECT 17.05 61.143 21.478 61.852 ;
        RECT 17.05 61.143 21.432 61.898 ;
        RECT 17.05 61.143 21.386 61.944 ;
        RECT 17.05 61.143 21.34 61.99 ;
        RECT 17.05 61.143 21.294 62.036 ;
        RECT 17.05 61.143 21.248 62.082 ;
        RECT 17.05 61.143 21.202 62.128 ;
        RECT 17.05 61.143 21.156 62.174 ;
        RECT 17.05 61.143 21.11 62.22 ;
        RECT 17.05 61.143 21.064 62.266 ;
        RECT 17.05 61.143 21.018 62.312 ;
        RECT 17.05 61.143 20.972 62.358 ;
        RECT 17.05 61.143 20.926 62.404 ;
        RECT 17.05 61.143 20.88 62.45 ;
        RECT 17.05 61.143 20.834 62.496 ;
        RECT 17.05 61.143 20.788 62.542 ;
        RECT 17.05 61.143 20.742 62.588 ;
        RECT 17.05 61.143 20.696 62.634 ;
        RECT 17.05 61.143 20.65 80 ;
        RECT 57.588 20.605 80 20.65 ;
        RECT 61.166 17.05 80 20.65 ;
        RECT 57.542 20.651 62.657 20.66 ;
        RECT 57.542 20.651 62.638 20.692 ;
        RECT 56.116 22.077 61.166 22.159 ;
        RECT 56.162 22.031 61.212 22.118 ;
        RECT 61.13 17.068 61.166 22.159 ;
        RECT 56.07 22.123 61.13 22.2 ;
        RECT 56.208 21.985 61.258 22.072 ;
        RECT 61.084 17.109 61.13 22.2 ;
        RECT 56.024 22.169 61.084 22.246 ;
        RECT 56.254 21.939 61.304 22.026 ;
        RECT 61.038 17.155 61.084 22.246 ;
        RECT 55.978 22.215 61.038 22.292 ;
        RECT 56.3 21.893 61.35 21.98 ;
        RECT 60.992 17.201 61.038 22.292 ;
        RECT 55.932 22.261 60.992 22.338 ;
        RECT 56.346 21.847 61.396 21.934 ;
        RECT 60.946 17.247 60.992 22.338 ;
        RECT 55.886 22.307 60.946 22.384 ;
        RECT 56.392 21.801 61.442 21.888 ;
        RECT 60.9 17.293 60.946 22.384 ;
        RECT 55.84 22.353 60.9 22.43 ;
        RECT 56.438 21.755 61.488 21.842 ;
        RECT 60.854 17.339 60.9 22.43 ;
        RECT 55.794 22.399 60.854 22.476 ;
        RECT 56.484 21.709 61.534 21.796 ;
        RECT 60.808 17.385 60.854 22.476 ;
        RECT 55.748 22.445 60.808 22.522 ;
        RECT 56.53 21.663 61.58 21.75 ;
        RECT 60.762 17.431 60.808 22.522 ;
        RECT 55.702 22.491 60.762 22.568 ;
        RECT 56.576 21.617 61.626 21.704 ;
        RECT 60.716 17.477 60.762 22.568 ;
        RECT 55.656 22.537 60.716 22.614 ;
        RECT 56.622 21.571 61.672 21.658 ;
        RECT 60.67 17.523 60.716 22.614 ;
        RECT 55.61 22.583 60.67 22.66 ;
        RECT 56.668 21.525 61.718 21.612 ;
        RECT 60.624 17.569 60.67 22.66 ;
        RECT 55.564 22.629 60.624 22.706 ;
        RECT 56.714 21.479 61.764 21.566 ;
        RECT 60.578 17.615 60.624 22.706 ;
        RECT 55.518 22.675 60.578 22.752 ;
        RECT 56.76 21.433 61.81 21.52 ;
        RECT 60.532 17.661 60.578 22.752 ;
        RECT 55.472 22.721 60.532 22.798 ;
        RECT 56.806 21.387 61.856 21.474 ;
        RECT 60.486 17.707 60.532 22.798 ;
        RECT 55.426 22.767 60.486 22.844 ;
        RECT 56.852 21.341 61.902 21.428 ;
        RECT 60.44 17.753 60.486 22.844 ;
        RECT 55.38 22.813 60.44 22.89 ;
        RECT 56.898 21.295 61.948 21.382 ;
        RECT 60.394 17.799 60.44 22.89 ;
        RECT 55.334 22.859 60.394 22.936 ;
        RECT 56.944 21.249 61.994 21.336 ;
        RECT 60.348 17.845 60.394 22.936 ;
        RECT 55.288 22.905 60.348 22.982 ;
        RECT 56.99 21.203 62.04 21.29 ;
        RECT 60.302 17.891 60.348 22.982 ;
        RECT 55.242 22.951 60.302 23.028 ;
        RECT 57.036 21.157 62.086 21.244 ;
        RECT 60.256 17.937 60.302 23.028 ;
        RECT 55.196 22.997 60.256 23.074 ;
        RECT 57.082 21.111 62.132 21.198 ;
        RECT 60.21 17.983 60.256 23.074 ;
        RECT 55.15 23.043 60.21 23.12 ;
        RECT 57.128 21.065 62.178 21.152 ;
        RECT 60.164 18.029 60.21 23.12 ;
        RECT 55.104 23.089 60.164 23.166 ;
        RECT 57.174 21.019 62.224 21.106 ;
        RECT 60.118 18.075 60.164 23.166 ;
        RECT 55.058 23.135 60.118 23.212 ;
        RECT 57.22 20.973 62.27 21.06 ;
        RECT 60.072 18.121 60.118 23.212 ;
        RECT 55.012 23.181 60.072 23.258 ;
        RECT 57.266 20.927 62.316 21.014 ;
        RECT 60.026 18.167 60.072 23.258 ;
        RECT 54.966 23.227 60.026 23.304 ;
        RECT 57.312 20.881 62.362 20.968 ;
        RECT 59.98 18.213 60.026 23.304 ;
        RECT 54.92 23.273 59.98 23.35 ;
        RECT 57.358 20.835 62.408 20.922 ;
        RECT 59.934 18.259 59.98 23.35 ;
        RECT 54.874 23.319 59.934 23.396 ;
        RECT 57.404 20.789 62.454 20.876 ;
        RECT 59.888 18.305 59.934 23.396 ;
        RECT 54.828 23.365 59.888 23.442 ;
        RECT 57.45 20.743 62.5 20.83 ;
        RECT 59.842 18.351 59.888 23.442 ;
        RECT 54.782 23.411 59.842 23.488 ;
        RECT 57.496 20.697 62.546 20.784 ;
        RECT 59.796 18.397 59.842 23.488 ;
        RECT 54.736 23.457 59.796 23.534 ;
        RECT 57.542 20.651 62.592 20.738 ;
        RECT 59.75 18.443 59.796 23.534 ;
        RECT 54.69 23.503 59.75 23.58 ;
        RECT 57.634 20.559 80 20.65 ;
        RECT 59.704 18.489 59.75 23.58 ;
        RECT 54.644 23.549 59.704 23.626 ;
        RECT 57.68 20.513 80 20.65 ;
        RECT 59.658 18.535 59.704 23.626 ;
        RECT 54.598 23.595 59.658 23.672 ;
        RECT 57.726 20.467 80 20.65 ;
        RECT 59.612 18.581 59.658 23.672 ;
        RECT 54.552 23.641 59.612 23.718 ;
        RECT 57.772 20.421 80 20.65 ;
        RECT 59.566 18.627 59.612 23.718 ;
        RECT 54.506 23.687 59.566 23.764 ;
        RECT 57.818 20.375 80 20.65 ;
        RECT 59.52 18.673 59.566 23.764 ;
        RECT 54.46 23.733 59.52 23.81 ;
        RECT 57.864 20.329 80 20.65 ;
        RECT 59.474 18.719 59.52 23.81 ;
        RECT 54.414 23.779 59.474 23.856 ;
        RECT 57.91 20.283 80 20.65 ;
        RECT 59.428 18.765 59.474 23.856 ;
        RECT 54.368 23.825 59.428 23.902 ;
        RECT 57.956 20.237 80 20.65 ;
        RECT 59.382 18.811 59.428 23.902 ;
        RECT 54.322 23.871 59.382 23.948 ;
        RECT 58.002 20.191 80 20.65 ;
        RECT 59.336 18.857 59.382 23.948 ;
        RECT 54.276 23.917 59.336 23.994 ;
        RECT 58.048 20.145 80 20.65 ;
        RECT 59.29 18.903 59.336 23.994 ;
        RECT 54.23 23.963 59.29 24.04 ;
        RECT 58.094 20.099 80 20.65 ;
        RECT 59.244 18.949 59.29 24.04 ;
        RECT 54.184 24.009 59.244 24.086 ;
        RECT 58.14 20.053 80 20.65 ;
        RECT 59.198 18.995 59.244 24.086 ;
        RECT 54.138 24.055 59.198 24.132 ;
        RECT 58.186 20.007 80 20.65 ;
        RECT 59.152 19.041 59.198 24.132 ;
        RECT 54.092 24.101 59.152 24.178 ;
        RECT 58.232 19.961 80 20.65 ;
        RECT 59.106 19.087 59.152 24.178 ;
        RECT 54.046 24.147 59.106 24.224 ;
        RECT 58.278 19.915 80 20.65 ;
        RECT 59.06 19.133 59.106 24.224 ;
        RECT 54 24.193 59.06 24.27 ;
        RECT 58.324 19.869 80 20.65 ;
        RECT 59.014 19.179 59.06 24.27 ;
        RECT 53.954 24.239 59.014 24.316 ;
        RECT 58.37 19.823 80 20.65 ;
        RECT 58.968 19.225 59.014 24.316 ;
        RECT 53.908 24.285 58.968 24.362 ;
        RECT 58.416 19.777 80 20.65 ;
        RECT 58.922 19.271 58.968 24.362 ;
        RECT 53.862 24.331 58.922 24.408 ;
        RECT 58.462 19.731 80 20.65 ;
        RECT 58.876 19.317 58.922 24.408 ;
        RECT 53.816 24.377 58.876 24.454 ;
        RECT 58.508 19.685 80 20.65 ;
        RECT 58.83 19.363 58.876 24.454 ;
        RECT 53.77 24.423 58.83 24.5 ;
        RECT 58.554 19.639 80 20.65 ;
        RECT 58.784 19.409 58.83 24.5 ;
        RECT 53.724 24.469 58.784 24.546 ;
        RECT 58.6 19.593 80 20.65 ;
        RECT 58.738 19.455 58.784 24.546 ;
        RECT 53.678 24.515 58.738 24.592 ;
        RECT 58.646 19.547 80 20.65 ;
        RECT 58.692 19.501 58.738 24.592 ;
        RECT 53.632 24.561 58.692 24.638 ;
        RECT 53.586 24.607 58.646 24.684 ;
        RECT 53.54 24.653 58.6 24.73 ;
        RECT 53.494 24.699 58.554 24.776 ;
        RECT 53.448 24.745 58.508 24.822 ;
        RECT 53.402 24.791 58.462 24.868 ;
        RECT 53.356 24.837 58.416 24.914 ;
        RECT 53.31 24.883 58.37 24.96 ;
        RECT 53.264 24.929 58.324 25.006 ;
        RECT 53.218 24.975 58.278 25.052 ;
        RECT 53.172 25.021 58.232 25.098 ;
        RECT 53.126 25.067 58.186 25.144 ;
        RECT 53.08 25.113 58.14 25.19 ;
        RECT 53.034 25.159 58.094 25.236 ;
        RECT 52.988 25.205 58.048 25.282 ;
        RECT 52.942 25.251 58.002 25.328 ;
        RECT 52.896 25.297 57.956 25.374 ;
        RECT 52.85 25.343 57.91 25.42 ;
        RECT 52.804 25.389 57.864 25.466 ;
        RECT 52.758 25.435 57.818 25.512 ;
        RECT 52.712 25.481 57.772 25.558 ;
        RECT 52.666 25.527 57.726 25.604 ;
        RECT 52.62 25.573 57.68 25.65 ;
        RECT 52.574 25.619 57.634 25.696 ;
        RECT 52.528 25.665 57.588 25.742 ;
        RECT 52.482 25.711 57.542 25.788 ;
        RECT 52.436 25.757 57.496 25.834 ;
        RECT 52.39 25.803 57.45 25.88 ;
        RECT 52.344 25.849 57.404 25.926 ;
        RECT 52.298 25.895 57.358 25.972 ;
        RECT 52.252 25.941 57.312 26.018 ;
        RECT 52.206 25.987 57.266 26.064 ;
        RECT 52.16 26.033 57.22 26.11 ;
        RECT 52.114 26.079 57.174 26.156 ;
        RECT 52.068 26.125 57.128 26.202 ;
        RECT 52.022 26.171 57.082 26.248 ;
        RECT 51.976 26.217 57.036 26.294 ;
        RECT 51.93 26.263 56.99 26.34 ;
        RECT 51.884 26.309 56.944 26.386 ;
        RECT 51.838 26.355 56.898 26.432 ;
        RECT 51.792 26.401 56.852 26.478 ;
        RECT 51.746 26.447 56.806 26.524 ;
        RECT 51.7 26.493 56.76 26.57 ;
        RECT 51.654 26.539 56.714 26.616 ;
        RECT 51.608 26.585 56.668 26.662 ;
        RECT 51.562 26.631 56.622 26.708 ;
        RECT 51.516 26.677 56.576 26.754 ;
        RECT 51.47 26.723 56.53 26.8 ;
        RECT 51.424 26.769 56.484 26.846 ;
        RECT 51.378 26.815 56.438 26.892 ;
        RECT 51.332 26.861 56.392 26.938 ;
        RECT 51.286 26.907 56.346 26.984 ;
        RECT 51.24 26.953 56.3 27.03 ;
        RECT 51.194 26.999 56.254 27.076 ;
        RECT 51.148 27.045 56.208 27.122 ;
        RECT 51.102 27.091 56.162 27.168 ;
        RECT 51.056 27.137 56.116 27.214 ;
        RECT 51.01 27.183 56.07 27.26 ;
        RECT 50.964 27.229 56.024 27.306 ;
        RECT 50.918 27.275 55.978 27.352 ;
        RECT 50.872 27.321 55.932 27.398 ;
        RECT 50.826 27.367 55.886 27.444 ;
        RECT 50.78 27.413 55.84 27.49 ;
        RECT 50.734 27.459 55.794 27.536 ;
        RECT 50.688 27.505 55.748 27.582 ;
        RECT 50.642 27.551 55.702 27.628 ;
        RECT 50.596 27.597 55.656 27.674 ;
        RECT 50.55 27.643 55.61 27.72 ;
        RECT 50.504 27.689 55.564 27.766 ;
        RECT 50.458 27.735 55.518 27.812 ;
        RECT 50.412 27.781 55.472 27.858 ;
        RECT 50.366 27.827 55.426 27.904 ;
        RECT 50.32 27.873 55.38 27.95 ;
        RECT 50.274 27.919 55.334 27.996 ;
        RECT 50.228 27.965 55.288 28.042 ;
        RECT 50.182 28.011 55.242 28.088 ;
        RECT 50.136 28.057 55.196 28.134 ;
        RECT 50.09 28.103 55.15 28.18 ;
        RECT 50.044 28.149 55.104 28.226 ;
        RECT 49.998 28.195 55.058 28.272 ;
        RECT 49.952 28.241 55.012 28.318 ;
        RECT 49.906 28.287 54.966 28.364 ;
        RECT 49.86 28.333 54.92 28.41 ;
        RECT 49.814 28.379 54.874 28.456 ;
        RECT 49.768 28.425 54.828 28.502 ;
        RECT 49.722 28.471 54.782 28.548 ;
        RECT 49.676 28.517 54.736 28.594 ;
        RECT 49.63 28.563 54.69 28.64 ;
        RECT 49.584 28.609 54.644 28.686 ;
        RECT 49.538 28.655 54.598 28.732 ;
        RECT 49.492 28.701 54.552 28.778 ;
        RECT 49.446 28.747 54.506 28.824 ;
        RECT 49.4 28.793 54.46 28.87 ;
        RECT 49.354 28.839 54.414 28.916 ;
        RECT 49.308 28.885 54.368 28.962 ;
        RECT 49.262 28.931 54.322 29.008 ;
        RECT 49.216 28.977 54.276 29.054 ;
        RECT 49.17 29.023 54.23 29.1 ;
        RECT 49.124 29.069 54.184 29.146 ;
        RECT 49.078 29.115 54.138 29.192 ;
        RECT 49.032 29.161 54.092 29.238 ;
        RECT 48.986 29.207 54.046 29.284 ;
        RECT 48.94 29.253 54 29.33 ;
        RECT 48.894 29.299 53.954 29.376 ;
        RECT 48.848 29.345 53.908 29.422 ;
        RECT 48.802 29.391 53.862 29.468 ;
        RECT 48.756 29.437 53.816 29.514 ;
        RECT 48.71 29.483 53.77 29.56 ;
        RECT 48.664 29.529 53.724 29.606 ;
        RECT 48.618 29.575 53.678 29.652 ;
        RECT 48.572 29.621 53.632 29.698 ;
        RECT 48.526 29.667 53.586 29.744 ;
        RECT 48.48 29.713 53.54 29.79 ;
        RECT 48.434 29.759 53.494 29.836 ;
        RECT 48.388 29.805 53.448 29.882 ;
        RECT 48.342 29.851 53.402 29.928 ;
        RECT 48.296 29.897 53.356 29.974 ;
        RECT 48.25 29.943 53.31 30.02 ;
        RECT 48.204 29.989 53.264 30.066 ;
        RECT 48.158 30.035 53.218 30.112 ;
        RECT 48.112 30.081 53.172 30.158 ;
        RECT 48.066 30.127 53.126 30.204 ;
        RECT 48.02 30.173 53.08 30.25 ;
        RECT 47.974 30.219 53.034 30.296 ;
        RECT 47.928 30.265 52.988 30.342 ;
        RECT 47.882 30.311 52.942 30.388 ;
        RECT 47.836 30.357 52.896 30.434 ;
        RECT 47.79 30.403 52.85 30.48 ;
        RECT 47.744 30.449 52.804 30.526 ;
        RECT 47.698 30.495 52.758 30.572 ;
        RECT 47.652 30.541 52.712 30.618 ;
        RECT 47.606 30.587 52.666 30.664 ;
        RECT 47.56 30.633 52.62 30.71 ;
        RECT 47.514 30.679 52.574 30.756 ;
        RECT 47.468 30.725 52.528 30.802 ;
        RECT 47.422 30.771 52.482 30.848 ;
        RECT 47.376 30.817 52.436 30.894 ;
        RECT 47.33 30.863 52.39 30.94 ;
        RECT 47.284 30.909 52.344 30.986 ;
        RECT 47.238 30.955 52.298 31.032 ;
        RECT 47.192 31.001 52.252 31.078 ;
        RECT 47.146 31.047 52.206 31.124 ;
        RECT 47.1 31.093 52.16 31.17 ;
        RECT 47.054 31.139 52.114 31.216 ;
        RECT 47.008 31.185 52.068 31.262 ;
        RECT 46.962 31.231 52.022 31.308 ;
        RECT 46.916 31.277 51.976 31.354 ;
        RECT 46.87 31.323 51.93 31.4 ;
        RECT 46.824 31.369 51.884 31.446 ;
        RECT 46.778 31.415 51.838 31.492 ;
        RECT 46.732 31.461 51.792 31.538 ;
        RECT 46.686 31.507 51.746 31.584 ;
        RECT 46.64 31.553 51.7 31.63 ;
        RECT 46.594 31.599 51.654 31.676 ;
        RECT 46.548 31.645 51.608 31.722 ;
        RECT 46.502 31.691 51.562 31.768 ;
        RECT 46.456 31.737 51.516 31.814 ;
        RECT 46.41 31.783 51.47 31.86 ;
        RECT 46.364 31.829 51.424 31.906 ;
        RECT 46.318 31.875 51.378 31.952 ;
        RECT 46.272 31.921 51.332 31.998 ;
        RECT 46.226 31.967 51.286 32.044 ;
        RECT 46.18 32.013 51.24 32.09 ;
        RECT 46.134 32.059 51.194 32.136 ;
        RECT 46.088 32.105 51.148 32.182 ;
        RECT 46.042 32.151 51.102 32.228 ;
        RECT 45.996 32.197 51.056 32.274 ;
        RECT 45.95 32.243 51.01 32.32 ;
        RECT 45.904 32.289 50.964 32.366 ;
        RECT 45.858 32.335 50.918 32.412 ;
        RECT 45.812 32.381 50.872 32.458 ;
        RECT 45.766 32.427 50.826 32.504 ;
        RECT 45.72 32.473 50.78 32.55 ;
        RECT 45.674 32.519 50.734 32.596 ;
        RECT 45.628 32.565 50.688 32.642 ;
        RECT 45.582 32.611 50.642 32.688 ;
        RECT 45.536 32.657 50.596 32.734 ;
        RECT 45.49 32.703 50.55 32.78 ;
        RECT 45.444 32.749 50.504 32.826 ;
        RECT 45.398 32.795 50.458 32.872 ;
        RECT 45.352 32.841 50.412 32.918 ;
        RECT 45.306 32.887 50.366 32.964 ;
        RECT 45.26 32.933 50.32 33.01 ;
        RECT 45.214 32.979 50.274 33.056 ;
        RECT 45.168 33.025 50.228 33.102 ;
        RECT 45.122 33.071 50.182 33.148 ;
        RECT 45.076 33.117 50.136 33.194 ;
        RECT 45.03 33.163 50.09 33.24 ;
        RECT 44.984 33.209 50.044 33.286 ;
        RECT 44.938 33.255 49.998 33.332 ;
        RECT 44.892 33.301 49.952 33.378 ;
        RECT 44.846 33.347 49.906 33.424 ;
        RECT 44.8 33.393 49.86 33.47 ;
        RECT 44.754 33.439 49.814 33.516 ;
        RECT 44.708 33.485 49.768 33.562 ;
        RECT 44.662 33.531 49.722 33.608 ;
        RECT 44.616 33.577 49.676 33.654 ;
        RECT 44.57 33.623 49.63 33.7 ;
        RECT 44.524 33.669 49.584 33.746 ;
        RECT 44.478 33.715 49.538 33.792 ;
        RECT 44.432 33.761 49.492 33.838 ;
        RECT 44.386 33.807 49.446 33.884 ;
        RECT 44.34 33.853 49.4 33.93 ;
        RECT 44.294 33.899 49.354 33.976 ;
        RECT 44.248 33.945 49.308 34.022 ;
        RECT 44.202 33.991 49.262 34.068 ;
        RECT 44.156 34.037 49.216 34.114 ;
        RECT 44.11 34.083 49.17 34.16 ;
        RECT 44.064 34.129 49.124 34.206 ;
        RECT 44.018 34.175 49.078 34.252 ;
        RECT 43.972 34.221 49.032 34.298 ;
        RECT 43.926 34.267 48.986 34.344 ;
        RECT 43.88 34.313 48.94 34.39 ;
        RECT 43.834 34.359 48.894 34.436 ;
        RECT 43.788 34.405 48.848 34.482 ;
        RECT 43.742 34.451 48.802 34.528 ;
        RECT 43.696 34.497 48.756 34.574 ;
        RECT 43.65 34.543 48.71 34.62 ;
        RECT 43.604 34.589 48.664 34.666 ;
        RECT 43.558 34.635 48.618 34.712 ;
        RECT 43.512 34.681 48.572 34.758 ;
        RECT 43.466 34.727 48.526 34.804 ;
        RECT 43.42 34.773 48.48 34.85 ;
        RECT 43.374 34.819 48.434 34.896 ;
        RECT 43.328 34.865 48.388 34.942 ;
        RECT 43.282 34.911 48.342 34.988 ;
        RECT 43.236 34.957 48.296 35.034 ;
        RECT 43.19 35.003 48.25 35.08 ;
        RECT 43.144 35.049 48.204 35.126 ;
        RECT 43.098 35.095 48.158 35.172 ;
        RECT 43.052 35.141 48.112 35.218 ;
        RECT 43.006 35.187 48.066 35.264 ;
        RECT 42.96 35.233 48.02 35.31 ;
        RECT 42.914 35.279 47.974 35.356 ;
        RECT 42.868 35.325 47.928 35.402 ;
        RECT 42.822 35.371 47.882 35.448 ;
        RECT 42.776 35.417 47.836 35.494 ;
        RECT 42.73 35.463 47.79 35.54 ;
        RECT 42.684 35.509 47.744 35.586 ;
        RECT 42.638 35.555 47.698 35.632 ;
        RECT 42.592 35.601 47.652 35.678 ;
        RECT 42.546 35.647 47.606 35.724 ;
        RECT 42.5 35.693 47.56 35.77 ;
        RECT 42.454 35.739 47.514 35.816 ;
        RECT 42.408 35.785 47.468 35.862 ;
        RECT 42.362 35.831 47.422 35.908 ;
        RECT 42.316 35.877 47.376 35.954 ;
        RECT 42.27 35.923 47.33 36 ;
        RECT 42.224 35.969 47.284 36.046 ;
        RECT 42.178 36.015 47.238 36.092 ;
        RECT 42.132 36.061 47.192 36.138 ;
        RECT 42.086 36.107 47.146 36.184 ;
        RECT 42.04 36.153 47.1 36.23 ;
        RECT 41.994 36.199 47.054 36.276 ;
        RECT 41.948 36.245 47.008 36.322 ;
        RECT 41.902 36.291 46.962 36.368 ;
        RECT 41.856 36.337 46.916 36.414 ;
        RECT 41.81 36.383 46.87 36.46 ;
        RECT 41.764 36.429 46.824 36.506 ;
        RECT 41.718 36.475 46.778 36.552 ;
        RECT 41.672 36.521 46.732 36.598 ;
        RECT 41.626 36.567 46.686 36.644 ;
        RECT 41.58 36.613 46.64 36.69 ;
        RECT 41.534 36.659 46.594 36.736 ;
        RECT 41.488 36.705 46.548 36.782 ;
        RECT 41.442 36.751 46.502 36.828 ;
        RECT 41.396 36.797 46.456 36.874 ;
        RECT 41.35 36.843 46.41 36.92 ;
        RECT 41.304 36.889 46.364 36.966 ;
        RECT 41.258 36.935 46.318 37.012 ;
        RECT 41.212 36.981 46.272 37.058 ;
        RECT 41.166 37.027 46.226 37.104 ;
        RECT 41.12 37.073 46.18 37.15 ;
        RECT 41.074 37.119 46.134 37.196 ;
        RECT 41.028 37.165 46.088 37.242 ;
        RECT 40.982 37.211 46.042 37.288 ;
        RECT 40.936 37.257 45.996 37.334 ;
        RECT 40.89 37.303 45.95 37.38 ;
        RECT 40.844 37.349 45.904 37.426 ;
        RECT 40.798 37.395 45.858 37.472 ;
        RECT 40.752 37.441 45.812 37.518 ;
        RECT 40.706 37.487 45.766 37.564 ;
        RECT 40.66 37.533 45.72 37.61 ;
        RECT 40.614 37.579 45.674 37.656 ;
        RECT 40.568 37.625 45.628 37.702 ;
        RECT 40.522 37.671 45.582 37.748 ;
        RECT 40.476 37.717 45.536 37.794 ;
        RECT 40.43 37.763 45.49 37.84 ;
        RECT 40.384 37.809 45.444 37.886 ;
        RECT 40.338 37.855 45.398 37.932 ;
        RECT 40.292 37.901 45.352 37.978 ;
        RECT 40.246 37.947 45.306 38.024 ;
        RECT 40.2 37.993 45.26 38.07 ;
        RECT 40.154 38.039 45.214 38.116 ;
        RECT 40.108 38.085 45.168 38.162 ;
        RECT 40.062 38.131 45.122 38.208 ;
        RECT 40.016 38.177 45.076 38.254 ;
        RECT 39.97 38.223 45.03 38.3 ;
        RECT 39.924 38.269 44.984 38.346 ;
        RECT 39.878 38.315 44.938 38.392 ;
        RECT 39.832 38.361 44.892 38.438 ;
        RECT 39.786 38.407 44.846 38.484 ;
        RECT 39.74 38.453 44.8 38.53 ;
        RECT 39.694 38.499 44.754 38.576 ;
        RECT 39.648 38.545 44.708 38.622 ;
        RECT 39.602 38.591 44.662 38.668 ;
        RECT 39.556 38.637 44.616 38.714 ;
        RECT 39.51 38.683 44.57 38.76 ;
        RECT 39.464 38.729 44.524 38.806 ;
        RECT 39.418 38.775 44.478 38.852 ;
        RECT 39.372 38.821 44.432 38.898 ;
        RECT 39.326 38.867 44.386 38.944 ;
        RECT 39.28 38.913 44.34 38.99 ;
        RECT 39.234 38.959 44.294 39.036 ;
        RECT 39.188 39.005 44.248 39.082 ;
        RECT 39.142 39.051 44.202 39.128 ;
        RECT 39.096 39.097 44.156 39.174 ;
        RECT 39.05 39.143 44.11 39.22 ;
        RECT 39.004 39.189 44.064 39.266 ;
        RECT 38.958 39.235 44.018 39.312 ;
        RECT 38.912 39.281 43.972 39.358 ;
        RECT 38.866 39.327 43.926 39.404 ;
        RECT 38.82 39.373 43.88 39.45 ;
        RECT 38.774 39.419 43.834 39.496 ;
        RECT 38.728 39.465 43.788 39.542 ;
        RECT 38.682 39.511 43.742 39.588 ;
        RECT 38.636 39.557 43.696 39.634 ;
        RECT 38.59 39.603 43.65 39.68 ;
        RECT 38.544 39.649 43.604 39.726 ;
        RECT 38.498 39.695 43.558 39.772 ;
        RECT 38.452 39.741 43.512 39.818 ;
        RECT 38.406 39.787 43.466 39.864 ;
        RECT 38.36 39.833 43.42 39.91 ;
        RECT 38.314 39.879 43.374 39.956 ;
        RECT 38.268 39.925 43.328 40.002 ;
        RECT 38.222 39.971 43.282 40.048 ;
        RECT 38.176 40.017 43.236 40.094 ;
        RECT 38.13 40.063 43.19 40.14 ;
        RECT 38.084 40.109 43.144 40.186 ;
        RECT 38.038 40.155 43.098 40.232 ;
        RECT 37.992 40.201 43.052 40.278 ;
        RECT 37.946 40.247 43.006 40.324 ;
        RECT 37.9 40.293 42.96 40.37 ;
        RECT 37.854 40.339 42.914 40.416 ;
        RECT 37.808 40.385 42.868 40.462 ;
        RECT 37.762 40.431 42.822 40.508 ;
        RECT 37.716 40.477 42.776 40.554 ;
        RECT 37.67 40.523 42.73 40.6 ;
        RECT 37.624 40.569 42.684 40.646 ;
        RECT 37.578 40.615 42.638 40.692 ;
        RECT 37.532 40.661 42.592 40.738 ;
        RECT 37.486 40.707 42.546 40.784 ;
        RECT 37.44 40.753 42.5 40.83 ;
        RECT 37.394 40.799 42.454 40.876 ;
        RECT 37.348 40.845 42.408 40.922 ;
        RECT 37.302 40.891 42.362 40.968 ;
        RECT 37.256 40.937 42.316 41.014 ;
        RECT 37.21 40.983 42.27 41.06 ;
        RECT 37.164 41.029 42.224 41.106 ;
        RECT 37.118 41.075 42.178 41.152 ;
        RECT 37.072 41.121 42.132 41.198 ;
        RECT 37.026 41.167 42.086 41.244 ;
        RECT 36.98 41.213 42.04 41.29 ;
        RECT 36.934 41.259 41.994 41.336 ;
        RECT 36.888 41.305 41.948 41.382 ;
        RECT 36.842 41.351 41.902 41.428 ;
        RECT 36.796 41.397 41.856 41.474 ;
        RECT 36.75 41.443 41.81 41.52 ;
        RECT 36.704 41.489 41.764 41.566 ;
        RECT 36.658 41.535 41.718 41.612 ;
        RECT 36.612 41.581 41.672 41.658 ;
        RECT 36.566 41.627 41.626 41.704 ;
        RECT 36.52 41.673 41.58 41.75 ;
        RECT 36.474 41.719 41.534 41.796 ;
        RECT 36.428 41.765 41.488 41.842 ;
        RECT 36.382 41.811 41.442 41.888 ;
        RECT 36.336 41.857 41.396 41.934 ;
        RECT 36.29 41.903 41.35 41.98 ;
        RECT 36.244 41.949 41.304 42.026 ;
        RECT 36.198 41.995 41.258 42.072 ;
        RECT 36.152 42.041 41.212 42.118 ;
        RECT 36.106 42.087 41.166 42.164 ;
        RECT 36.06 42.133 41.12 42.21 ;
        RECT 36.014 42.179 41.074 42.256 ;
        RECT 35.968 42.225 41.028 42.302 ;
        RECT 35.922 42.271 40.982 42.348 ;
        RECT 35.876 42.317 40.936 42.394 ;
        RECT 35.83 42.363 40.89 42.44 ;
        RECT 35.784 42.409 40.844 42.486 ;
        RECT 35.738 42.455 40.798 42.532 ;
        RECT 35.692 42.501 40.752 42.578 ;
        RECT 35.646 42.547 40.706 42.624 ;
        RECT 35.6 42.593 40.66 42.67 ;
        RECT 35.554 42.639 40.614 42.716 ;
        RECT 35.508 42.685 40.568 42.762 ;
        RECT 35.462 42.731 40.522 42.808 ;
        RECT 35.416 42.777 40.476 42.854 ;
        RECT 35.37 42.823 40.43 42.9 ;
        RECT 35.324 42.869 40.384 42.946 ;
        RECT 35.278 42.915 40.338 42.992 ;
        RECT 35.232 42.961 40.292 43.038 ;
        RECT 35.186 43.007 40.246 43.084 ;
        RECT 35.14 43.053 40.2 43.13 ;
        RECT 35.094 43.099 40.154 43.176 ;
        RECT 35.048 43.145 40.108 43.222 ;
        RECT 35.002 43.191 40.062 43.268 ;
        RECT 34.956 43.237 40.016 43.314 ;
        RECT 34.91 43.283 39.97 43.36 ;
        RECT 34.864 43.329 39.924 43.406 ;
        RECT 34.818 43.375 39.878 43.452 ;
        RECT 34.772 43.421 39.832 43.498 ;
        RECT 34.726 43.467 39.786 43.544 ;
        RECT 34.68 43.513 39.74 43.59 ;
        RECT 34.634 43.559 39.694 43.636 ;
        RECT 34.588 43.605 39.648 43.682 ;
        RECT 34.542 43.651 39.602 43.728 ;
        RECT 34.496 43.697 39.556 43.774 ;
        RECT 34.45 43.743 39.51 43.82 ;
        RECT 34.404 43.789 39.464 43.866 ;
        RECT 34.358 43.835 39.418 43.912 ;
        RECT 34.312 43.881 39.372 43.958 ;
        RECT 34.266 43.927 39.326 44.004 ;
        RECT 34.22 43.973 39.28 44.05 ;
        RECT 34.174 44.019 39.234 44.096 ;
        RECT 34.128 44.065 39.188 44.142 ;
        RECT 34.082 44.111 39.142 44.188 ;
        RECT 34.036 44.157 39.096 44.234 ;
        RECT 33.99 44.203 39.05 44.28 ;
        RECT 33.944 44.249 39.004 44.326 ;
        RECT 33.898 44.295 38.958 44.372 ;
        RECT 33.852 44.341 38.912 44.418 ;
        RECT 33.806 44.387 38.866 44.464 ;
        RECT 33.76 44.433 38.82 44.51 ;
        RECT 33.714 44.479 38.774 44.556 ;
        RECT 33.668 44.525 38.728 44.602 ;
        RECT 33.622 44.571 38.682 44.648 ;
        RECT 33.576 44.617 38.636 44.694 ;
        RECT 33.53 44.663 38.59 44.74 ;
        RECT 33.484 44.709 38.544 44.786 ;
        RECT 33.438 44.755 38.498 44.832 ;
        RECT 33.392 44.801 38.452 44.878 ;
        RECT 33.346 44.847 38.406 44.924 ;
        RECT 33.3 44.893 38.36 44.97 ;
        RECT 33.254 44.939 38.314 45.016 ;
        RECT 33.208 44.985 38.268 45.062 ;
        RECT 33.162 45.031 38.222 45.108 ;
        RECT 33.116 45.077 38.176 45.154 ;
        RECT 33.07 45.123 38.13 45.2 ;
        RECT 33.024 45.169 38.084 45.246 ;
        RECT 32.978 45.215 38.038 45.292 ;
        RECT 32.932 45.261 37.992 45.338 ;
        RECT 32.886 45.307 37.946 45.384 ;
        RECT 32.84 45.353 37.9 45.43 ;
        RECT 32.794 45.399 37.854 45.476 ;
        RECT 32.748 45.445 37.808 45.522 ;
        RECT 32.702 45.491 37.762 45.568 ;
        RECT 32.656 45.537 37.716 45.614 ;
        RECT 32.61 45.583 37.67 45.66 ;
        RECT 32.564 45.629 37.624 45.706 ;
        RECT 32.518 45.675 37.578 45.752 ;
        RECT 32.472 45.721 37.532 45.798 ;
        RECT 32.426 45.767 37.486 45.844 ;
        RECT 32.38 45.813 37.44 45.89 ;
        RECT 32.334 45.859 37.394 45.936 ;
        RECT 32.288 45.905 37.348 45.982 ;
        RECT 32.242 45.951 37.302 46.028 ;
        RECT 32.196 45.997 37.256 46.074 ;
        RECT 32.15 46.043 37.21 46.12 ;
        RECT 32.104 46.089 37.164 46.166 ;
        RECT 32.058 46.135 37.118 46.212 ;
        RECT 32.012 46.181 37.072 46.258 ;
        RECT 31.966 46.227 37.026 46.304 ;
        RECT 31.92 46.273 36.98 46.35 ;
        RECT 31.874 46.319 36.934 46.396 ;
        RECT 31.828 46.365 36.888 46.442 ;
        RECT 31.782 46.411 36.842 46.488 ;
        RECT 31.736 46.457 36.796 46.534 ;
        RECT 31.69 46.503 36.75 46.58 ;
        RECT 31.644 46.549 36.704 46.626 ;
        RECT 31.598 46.595 36.658 46.672 ;
        RECT 31.552 46.641 36.612 46.718 ;
        RECT 31.506 46.687 36.566 46.764 ;
        RECT 31.46 46.733 36.52 46.81 ;
        RECT 31.414 46.779 36.474 46.856 ;
        RECT 31.368 46.825 36.428 46.902 ;
        RECT 31.322 46.871 36.382 46.948 ;
        RECT 31.276 46.917 36.336 46.994 ;
        RECT 31.23 46.963 36.29 47.04 ;
        RECT 31.184 47.009 36.244 47.086 ;
        RECT 31.138 47.055 36.198 47.132 ;
        RECT 31.092 47.101 36.152 47.178 ;
        RECT 31.046 47.147 36.106 47.224 ;
        RECT 31 47.193 36.06 47.27 ;
        RECT 30.954 47.239 36.014 47.316 ;
        RECT 30.908 47.285 35.968 47.362 ;
        RECT 30.862 47.331 35.922 47.408 ;
        RECT 30.816 47.377 35.876 47.454 ;
        RECT 30.77 47.423 35.83 47.5 ;
        RECT 30.724 47.469 35.784 47.546 ;
        RECT 30.678 47.515 35.738 47.592 ;
        RECT 30.632 47.561 35.692 47.638 ;
        RECT 30.586 47.607 35.646 47.684 ;
        RECT 30.54 47.653 35.6 47.73 ;
        RECT 30.494 47.699 35.554 47.776 ;
        RECT 30.448 47.745 35.508 47.822 ;
        RECT 30.402 47.791 35.462 47.868 ;
        RECT 30.356 47.837 35.416 47.914 ;
        RECT 30.31 47.883 35.37 47.96 ;
        RECT 30.264 47.929 35.324 48.006 ;
        RECT 30.218 47.975 35.278 48.052 ;
        RECT 30.172 48.021 35.232 48.098 ;
        RECT 30.126 48.067 35.186 48.144 ;
        RECT 30.08 48.113 35.14 48.19 ;
        RECT 30.034 48.159 35.094 48.236 ;
        RECT 29.988 48.205 35.048 48.282 ;
        RECT 29.942 48.251 35.002 48.328 ;
        RECT 29.896 48.297 34.956 48.374 ;
        RECT 29.85 48.343 34.91 48.42 ;
        RECT 29.804 48.389 34.864 48.466 ;
        RECT 29.758 48.435 34.818 48.512 ;
        RECT 29.712 48.481 34.772 48.558 ;
        RECT 29.666 48.527 34.726 48.604 ;
        RECT 29.62 48.573 34.68 48.65 ;
        RECT 29.574 48.619 34.634 48.696 ;
        RECT 29.528 48.665 34.588 48.742 ;
        RECT 29.482 48.711 34.542 48.788 ;
        RECT 29.436 48.757 34.496 48.834 ;
        RECT 29.39 48.803 34.45 48.88 ;
        RECT 29.344 48.849 34.404 48.926 ;
        RECT 29.298 48.895 34.358 48.972 ;
        RECT 29.252 48.941 34.312 49.018 ;
        RECT 29.206 48.987 34.266 49.064 ;
        RECT 29.16 49.033 34.22 49.11 ;
        RECT 29.114 49.079 34.174 49.156 ;
        RECT 29.068 49.125 34.128 49.202 ;
        RECT 29.022 49.171 34.082 49.248 ;
        RECT 28.976 49.217 34.036 49.294 ;
        RECT 28.93 49.263 33.99 49.34 ;
        RECT 28.884 49.309 33.944 49.386 ;
        RECT 28.838 49.355 33.898 49.432 ;
        RECT 28.792 49.401 33.852 49.478 ;
        RECT 28.746 49.447 33.806 49.524 ;
        RECT 28.7 49.493 33.76 49.57 ;
        RECT 28.654 49.539 33.714 49.616 ;
        RECT 28.608 49.585 33.668 49.662 ;
        RECT 28.562 49.631 33.622 49.708 ;
        RECT 28.516 49.677 33.576 49.754 ;
        RECT 28.47 49.723 33.53 49.8 ;
        RECT 28.424 49.769 33.484 49.846 ;
        RECT 28.378 49.815 33.438 49.892 ;
        RECT 28.332 49.861 33.392 49.938 ;
        RECT 28.286 49.907 33.346 49.984 ;
        RECT 28.24 49.953 33.3 50.03 ;
        RECT 28.194 49.999 33.254 50.076 ;
        RECT 28.148 50.045 33.208 50.122 ;
        RECT 28.102 50.091 33.162 50.168 ;
        RECT 28.056 50.137 33.116 50.214 ;
        RECT 28.01 50.183 33.07 50.26 ;
        RECT 27.964 50.229 33.024 50.306 ;
        RECT 27.918 50.275 32.978 50.352 ;
        RECT 27.872 50.321 32.932 50.398 ;
        RECT 27.826 50.367 32.886 50.444 ;
        RECT 27.78 50.413 32.84 50.49 ;
        RECT 27.734 50.459 32.794 50.536 ;
        RECT 27.688 50.505 32.748 50.582 ;
        RECT 27.642 50.551 32.702 50.628 ;
        RECT 27.596 50.597 32.656 50.674 ;
        RECT 27.55 50.643 32.61 50.72 ;
        RECT 27.504 50.689 32.564 50.766 ;
        RECT 27.458 50.735 32.518 50.812 ;
        RECT 27.412 50.781 32.472 50.858 ;
        RECT 27.366 50.827 32.426 50.904 ;
        RECT 27.32 50.873 32.38 50.95 ;
        RECT 27.274 50.919 32.334 50.996 ;
        RECT 27.228 50.965 32.288 51.042 ;
        RECT 27.182 51.011 32.242 51.088 ;
        RECT 27.136 51.057 32.196 51.134 ;
        RECT 27.09 51.103 32.15 51.18 ;
        RECT 27.044 51.149 32.104 51.226 ;
        RECT 26.998 51.195 32.058 51.272 ;
        RECT 26.952 51.241 32.012 51.318 ;
        RECT 26.906 51.287 31.966 51.364 ;
        RECT 26.86 51.333 31.92 51.41 ;
        RECT 26.814 51.379 31.874 51.456 ;
        RECT 26.768 51.425 31.828 51.502 ;
        RECT 26.722 51.471 31.782 51.548 ;
        RECT 26.676 51.517 31.736 51.594 ;
        RECT 26.63 51.563 31.69 51.64 ;
        RECT 26.584 51.609 31.644 51.686 ;
        RECT 26.538 51.655 31.598 51.732 ;
        RECT 26.492 51.701 31.552 51.778 ;
        RECT 26.446 51.747 31.506 51.824 ;
        RECT 26.4 51.793 31.46 51.87 ;
        RECT 26.354 51.839 31.414 51.916 ;
        RECT 26.308 51.885 31.368 51.962 ;
        RECT 26.262 51.931 31.322 52.008 ;
        RECT 26.216 51.977 31.276 52.054 ;
        RECT 26.17 52.023 31.23 52.1 ;
        RECT 26.124 52.069 31.184 52.146 ;
        RECT 26.078 52.115 31.138 52.192 ;
        RECT 26.032 52.161 31.092 52.238 ;
        RECT 25.986 52.207 31.046 52.284 ;
        RECT 25.94 52.253 31 52.33 ;
        RECT 25.894 52.299 30.954 52.376 ;
        RECT 25.848 52.345 30.908 52.422 ;
        RECT 25.802 52.391 30.862 52.468 ;
        RECT 25.756 52.437 30.816 52.514 ;
        RECT 25.71 52.483 30.77 52.56 ;
        RECT 25.664 52.529 30.724 52.606 ;
        RECT 25.618 52.575 30.678 52.652 ;
        RECT 25.572 52.621 30.632 52.698 ;
        RECT 25.526 52.667 30.586 52.744 ;
        RECT 25.48 52.713 30.54 52.79 ;
        RECT 25.434 52.759 30.494 52.836 ;
        RECT 25.388 52.805 30.448 52.882 ;
        RECT 25.342 52.851 30.402 52.928 ;
        RECT 25.296 52.897 30.356 52.974 ;
        RECT 25.25 52.943 30.31 53.02 ;
        RECT 25.204 52.989 30.264 53.066 ;
        RECT 25.158 53.035 30.218 53.112 ;
        RECT 25.112 53.081 30.172 53.158 ;
        RECT 25.066 53.127 30.126 53.204 ;
        RECT 25.02 53.173 30.08 53.25 ;
        RECT 24.974 53.219 30.034 53.296 ;
        RECT 24.928 53.265 29.988 53.342 ;
        RECT 24.882 53.311 29.942 53.388 ;
        RECT 24.836 53.357 29.896 53.434 ;
        RECT 24.79 53.403 29.85 53.48 ;
        RECT 24.744 53.449 29.804 53.526 ;
        RECT 24.698 53.495 29.758 53.572 ;
        RECT 24.652 53.541 29.712 53.618 ;
        RECT 24.606 53.587 29.666 53.664 ;
        RECT 24.56 53.633 29.62 53.71 ;
        RECT 24.514 53.679 29.574 53.756 ;
        RECT 24.468 53.725 29.528 53.802 ;
        RECT 24.422 53.771 29.482 53.848 ;
        RECT 24.376 53.817 29.436 53.894 ;
        RECT 24.33 53.863 29.39 53.94 ;
        RECT 24.284 53.909 29.344 53.986 ;
        RECT 24.238 53.955 29.298 54.032 ;
        RECT 24.192 54.001 29.252 54.078 ;
        RECT 24.146 54.047 29.206 54.124 ;
        RECT 24.1 54.093 29.16 54.17 ;
        RECT 24.054 54.139 29.114 54.216 ;
        RECT 24.008 54.185 29.068 54.262 ;
        RECT 23.962 54.231 29.022 54.308 ;
        RECT 23.916 54.277 28.976 54.354 ;
        RECT 23.87 54.323 28.93 54.4 ;
        RECT 23.824 54.369 28.884 54.446 ;
        RECT 23.778 54.415 28.838 54.492 ;
        RECT 23.732 54.461 28.792 54.538 ;
        RECT 23.686 54.507 28.746 54.584 ;
        RECT 23.64 54.553 28.7 54.63 ;
        RECT 23.594 54.599 28.654 54.676 ;
        RECT 23.548 54.645 28.608 54.722 ;
        RECT 23.502 54.691 28.562 54.768 ;
        RECT 23.456 54.737 28.516 54.814 ;
        RECT 23.41 54.783 28.47 54.86 ;
        RECT 23.364 54.829 28.424 54.906 ;
        RECT 23.318 54.875 28.378 54.952 ;
        RECT 23.272 54.921 28.332 54.998 ;
        RECT 23.226 54.967 28.286 55.044 ;
        RECT 23.18 55.013 28.24 55.09 ;
        RECT 23.134 55.059 28.194 55.136 ;
        RECT 23.088 55.105 28.148 55.182 ;
        RECT 23.042 55.151 28.102 55.228 ;
        RECT 22.996 55.197 28.056 55.274 ;
        RECT 22.95 55.243 28.01 55.32 ;
        RECT 22.904 55.289 27.964 55.366 ;
        RECT 22.858 55.335 27.918 55.412 ;
        RECT 22.812 55.381 27.872 55.458 ;
        RECT 22.766 55.427 27.826 55.504 ;
        RECT 22.72 55.473 27.78 55.55 ;
        RECT 22.674 55.519 27.734 55.596 ;
        RECT 22.628 55.565 27.688 55.642 ;
        RECT 22.582 55.611 27.642 55.688 ;
    END
    PORT
      LAYER IB ;
        RECT 66.206 45.25 80 48.85 ;
        RECT 62.604 48.829 67.697 48.86 ;
        RECT 61.132 50.301 66.206 50.348 ;
        RECT 61.178 50.255 66.252 50.318 ;
        RECT 66.192 45.257 66.206 50.348 ;
        RECT 61.224 50.209 66.298 50.272 ;
        RECT 66.146 45.287 66.192 50.378 ;
        RECT 61.086 50.347 66.146 50.424 ;
        RECT 61.27 50.163 66.344 50.226 ;
        RECT 66.1 45.333 66.146 50.424 ;
        RECT 61.04 50.393 66.1 50.47 ;
        RECT 61.316 50.117 66.39 50.18 ;
        RECT 66.054 45.379 66.1 50.47 ;
        RECT 60.994 50.439 66.054 50.516 ;
        RECT 61.362 50.071 66.436 50.134 ;
        RECT 66.008 45.425 66.054 50.516 ;
        RECT 60.948 50.485 66.008 50.562 ;
        RECT 61.408 50.025 66.482 50.088 ;
        RECT 65.962 45.471 66.008 50.562 ;
        RECT 60.902 50.531 65.962 50.608 ;
        RECT 61.454 49.979 66.528 50.042 ;
        RECT 65.916 45.517 65.962 50.608 ;
        RECT 60.856 50.577 65.916 50.654 ;
        RECT 61.5 49.933 66.574 49.996 ;
        RECT 65.87 45.563 65.916 50.654 ;
        RECT 60.81 50.623 65.87 50.7 ;
        RECT 61.546 49.887 66.62 49.95 ;
        RECT 65.824 45.609 65.87 50.7 ;
        RECT 60.764 50.669 65.824 50.746 ;
        RECT 61.592 49.841 66.666 49.904 ;
        RECT 65.778 45.655 65.824 50.746 ;
        RECT 60.718 50.715 65.778 50.792 ;
        RECT 61.638 49.795 66.712 49.858 ;
        RECT 65.732 45.701 65.778 50.792 ;
        RECT 60.672 50.761 65.732 50.838 ;
        RECT 61.684 49.749 66.758 49.812 ;
        RECT 65.686 45.747 65.732 50.838 ;
        RECT 60.626 50.807 65.686 50.884 ;
        RECT 61.73 49.703 66.804 49.766 ;
        RECT 65.64 45.793 65.686 50.884 ;
        RECT 60.58 50.853 65.64 50.93 ;
        RECT 61.776 49.657 66.85 49.72 ;
        RECT 65.594 45.839 65.64 50.93 ;
        RECT 60.534 50.899 65.594 50.976 ;
        RECT 61.822 49.611 66.896 49.674 ;
        RECT 65.548 45.885 65.594 50.976 ;
        RECT 60.488 50.945 65.548 51.022 ;
        RECT 61.868 49.565 66.942 49.628 ;
        RECT 65.502 45.931 65.548 51.022 ;
        RECT 60.442 50.991 65.502 51.068 ;
        RECT 61.914 49.519 66.988 49.582 ;
        RECT 65.456 45.977 65.502 51.068 ;
        RECT 60.396 51.037 65.456 51.114 ;
        RECT 61.96 49.473 67.034 49.536 ;
        RECT 65.41 46.023 65.456 51.114 ;
        RECT 60.35 51.083 65.41 51.16 ;
        RECT 62.006 49.427 67.08 49.49 ;
        RECT 65.364 46.069 65.41 51.16 ;
        RECT 60.304 51.129 65.364 51.206 ;
        RECT 62.052 49.381 67.126 49.444 ;
        RECT 65.318 46.115 65.364 51.206 ;
        RECT 60.258 51.175 65.318 51.252 ;
        RECT 62.098 49.335 67.172 49.398 ;
        RECT 65.272 46.161 65.318 51.252 ;
        RECT 60.212 51.221 65.272 51.298 ;
        RECT 62.144 49.289 67.218 49.352 ;
        RECT 65.226 46.207 65.272 51.298 ;
        RECT 60.166 51.267 65.226 51.344 ;
        RECT 62.19 49.243 67.264 49.306 ;
        RECT 65.18 46.253 65.226 51.344 ;
        RECT 60.12 51.313 65.18 51.39 ;
        RECT 62.236 49.197 67.31 49.26 ;
        RECT 65.134 46.299 65.18 51.39 ;
        RECT 60.074 51.359 65.134 51.436 ;
        RECT 62.282 49.151 67.356 49.214 ;
        RECT 65.088 46.345 65.134 51.436 ;
        RECT 60.028 51.405 65.088 51.482 ;
        RECT 62.328 49.105 67.402 49.168 ;
        RECT 65.042 46.391 65.088 51.482 ;
        RECT 59.982 51.451 65.042 51.528 ;
        RECT 62.374 49.059 67.448 49.122 ;
        RECT 64.996 46.437 65.042 51.528 ;
        RECT 59.936 51.497 64.996 51.574 ;
        RECT 62.42 49.013 67.494 49.076 ;
        RECT 64.95 46.483 64.996 51.574 ;
        RECT 59.89 51.543 64.95 51.62 ;
        RECT 62.466 48.967 67.54 49.03 ;
        RECT 64.904 46.529 64.95 51.62 ;
        RECT 59.844 51.589 64.904 51.666 ;
        RECT 62.512 48.921 67.586 48.984 ;
        RECT 64.858 46.575 64.904 51.666 ;
        RECT 59.798 51.635 64.858 51.712 ;
        RECT 62.558 48.875 67.632 48.938 ;
        RECT 64.812 46.621 64.858 51.712 ;
        RECT 59.752 51.681 64.812 51.758 ;
        RECT 62.604 48.829 67.678 48.892 ;
        RECT 64.766 46.667 64.812 51.758 ;
        RECT 59.706 51.727 64.766 51.804 ;
        RECT 62.65 48.783 80 48.85 ;
        RECT 64.72 46.713 64.766 51.804 ;
        RECT 59.66 51.773 64.72 51.85 ;
        RECT 62.696 48.737 80 48.85 ;
        RECT 64.674 46.759 64.72 51.85 ;
        RECT 59.614 51.819 64.674 51.896 ;
        RECT 62.742 48.691 80 48.85 ;
        RECT 64.628 46.805 64.674 51.896 ;
        RECT 59.568 51.865 64.628 51.942 ;
        RECT 62.788 48.645 80 48.85 ;
        RECT 64.582 46.851 64.628 51.942 ;
        RECT 59.522 51.911 64.582 51.988 ;
        RECT 62.834 48.599 80 48.85 ;
        RECT 64.536 46.897 64.582 51.988 ;
        RECT 59.476 51.957 64.536 52.034 ;
        RECT 62.88 48.553 80 48.85 ;
        RECT 64.49 46.943 64.536 52.034 ;
        RECT 59.43 52.003 64.49 52.08 ;
        RECT 62.926 48.507 80 48.85 ;
        RECT 64.444 46.989 64.49 52.08 ;
        RECT 59.384 52.049 64.444 52.126 ;
        RECT 62.972 48.461 80 48.85 ;
        RECT 64.398 47.035 64.444 52.126 ;
        RECT 59.338 52.095 64.398 52.172 ;
        RECT 63.018 48.415 80 48.85 ;
        RECT 64.352 47.081 64.398 52.172 ;
        RECT 59.292 52.141 64.352 52.218 ;
        RECT 63.064 48.369 80 48.85 ;
        RECT 64.306 47.127 64.352 52.218 ;
        RECT 59.246 52.187 64.306 52.264 ;
        RECT 63.11 48.323 80 48.85 ;
        RECT 64.26 47.173 64.306 52.264 ;
        RECT 59.2 52.233 64.26 52.31 ;
        RECT 63.156 48.277 80 48.85 ;
        RECT 64.214 47.219 64.26 52.31 ;
        RECT 59.154 52.279 64.214 52.356 ;
        RECT 63.202 48.231 80 48.85 ;
        RECT 64.168 47.265 64.214 52.356 ;
        RECT 59.108 52.325 64.168 52.402 ;
        RECT 63.248 48.185 80 48.85 ;
        RECT 64.122 47.311 64.168 52.402 ;
        RECT 59.062 52.371 64.122 52.448 ;
        RECT 63.294 48.139 80 48.85 ;
        RECT 64.076 47.357 64.122 52.448 ;
        RECT 59.016 52.417 64.076 52.494 ;
        RECT 63.34 48.093 80 48.85 ;
        RECT 64.03 47.403 64.076 52.494 ;
        RECT 58.97 52.463 64.03 52.54 ;
        RECT 63.386 48.047 80 48.85 ;
        RECT 63.984 47.449 64.03 52.54 ;
        RECT 58.924 52.509 63.984 52.586 ;
        RECT 63.432 48.001 80 48.85 ;
        RECT 63.938 47.495 63.984 52.586 ;
        RECT 58.878 52.555 63.938 52.632 ;
        RECT 63.478 47.955 80 48.85 ;
        RECT 63.892 47.541 63.938 52.632 ;
        RECT 58.832 52.601 63.892 52.678 ;
        RECT 63.524 47.909 80 48.85 ;
        RECT 63.846 47.587 63.892 52.678 ;
        RECT 58.786 52.647 63.846 52.724 ;
        RECT 63.57 47.863 80 48.85 ;
        RECT 63.8 47.633 63.846 52.724 ;
        RECT 58.74 52.693 63.8 52.77 ;
        RECT 63.616 47.817 80 48.85 ;
        RECT 63.754 47.679 63.8 52.77 ;
        RECT 58.694 52.739 63.754 52.816 ;
        RECT 63.662 47.771 80 48.85 ;
        RECT 63.708 47.725 63.754 52.816 ;
        RECT 58.648 52.785 63.708 52.862 ;
        RECT 58.602 52.831 63.662 52.908 ;
        RECT 58.556 52.877 63.616 52.954 ;
        RECT 58.51 52.923 63.57 53 ;
        RECT 58.464 52.969 63.524 53.046 ;
        RECT 58.418 53.015 63.478 53.092 ;
        RECT 58.372 53.061 63.432 53.138 ;
        RECT 58.326 53.107 63.386 53.184 ;
        RECT 58.28 53.153 63.34 53.23 ;
        RECT 58.234 53.199 63.294 53.276 ;
        RECT 58.188 53.245 63.248 53.322 ;
        RECT 58.142 53.291 63.202 53.368 ;
        RECT 58.096 53.337 63.156 53.414 ;
        RECT 58.05 53.383 63.11 53.46 ;
        RECT 58.004 53.429 63.064 53.506 ;
        RECT 57.958 53.475 63.018 53.552 ;
        RECT 57.912 53.521 62.972 53.598 ;
        RECT 57.866 53.567 62.926 53.644 ;
        RECT 57.82 53.613 62.88 53.69 ;
        RECT 57.774 53.659 62.834 53.736 ;
        RECT 57.728 53.705 62.788 53.782 ;
        RECT 57.682 53.751 62.742 53.828 ;
        RECT 57.636 53.797 62.696 53.874 ;
        RECT 57.59 53.843 62.65 53.92 ;
        RECT 57.544 53.889 62.604 53.966 ;
        RECT 57.498 53.935 62.558 54.012 ;
        RECT 57.452 53.981 62.512 54.058 ;
        RECT 57.406 54.027 62.466 54.104 ;
        RECT 57.36 54.073 62.42 54.15 ;
        RECT 57.314 54.119 62.374 54.196 ;
        RECT 57.268 54.165 62.328 54.242 ;
        RECT 57.222 54.211 62.282 54.288 ;
        RECT 57.176 54.257 62.236 54.334 ;
        RECT 57.13 54.303 62.19 54.38 ;
        RECT 57.084 54.349 62.144 54.426 ;
        RECT 57.038 54.395 62.098 54.472 ;
        RECT 56.992 54.441 62.052 54.518 ;
        RECT 56.946 54.487 62.006 54.564 ;
        RECT 56.9 54.533 61.96 54.61 ;
        RECT 56.854 54.579 61.914 54.656 ;
        RECT 56.808 54.625 61.868 54.702 ;
        RECT 56.762 54.671 61.822 54.748 ;
        RECT 56.716 54.717 61.776 54.794 ;
        RECT 56.67 54.763 61.73 54.84 ;
        RECT 56.624 54.809 61.684 54.886 ;
        RECT 56.578 54.855 61.638 54.932 ;
        RECT 56.532 54.901 61.592 54.978 ;
        RECT 56.486 54.947 61.546 55.024 ;
        RECT 56.44 54.993 61.5 55.07 ;
        RECT 56.394 55.039 61.454 55.116 ;
        RECT 56.348 55.085 61.408 55.162 ;
        RECT 56.302 55.131 61.362 55.208 ;
        RECT 56.256 55.177 61.316 55.254 ;
        RECT 56.21 55.223 61.27 55.3 ;
        RECT 56.164 55.269 61.224 55.346 ;
        RECT 56.118 55.315 61.178 55.392 ;
        RECT 56.072 55.361 61.132 55.438 ;
        RECT 56.026 55.407 61.086 55.484 ;
        RECT 55.98 55.453 61.04 55.53 ;
        RECT 55.934 55.499 60.994 55.576 ;
        RECT 55.888 55.545 60.948 55.622 ;
        RECT 55.842 55.591 60.902 55.668 ;
        RECT 55.796 55.637 60.856 55.714 ;
        RECT 55.75 55.683 60.81 55.76 ;
        RECT 55.704 55.729 60.764 55.806 ;
        RECT 55.658 55.775 60.718 55.852 ;
        RECT 55.612 55.821 60.672 55.898 ;
        RECT 55.566 55.867 60.626 55.944 ;
        RECT 55.52 55.913 60.58 55.99 ;
        RECT 55.474 55.959 60.534 56.036 ;
        RECT 55.428 56.005 60.488 56.082 ;
        RECT 55.382 56.051 60.442 56.128 ;
        RECT 55.336 56.097 60.396 56.174 ;
        RECT 55.29 56.143 60.35 56.22 ;
        RECT 55.244 56.189 60.304 56.266 ;
        RECT 55.198 56.235 60.258 56.312 ;
        RECT 55.152 56.281 60.212 56.358 ;
        RECT 55.106 56.327 60.166 56.404 ;
        RECT 55.06 56.373 60.12 56.45 ;
        RECT 55.014 56.419 60.074 56.496 ;
        RECT 54.968 56.465 60.028 56.542 ;
        RECT 54.922 56.511 59.982 56.588 ;
        RECT 54.876 56.557 59.936 56.634 ;
        RECT 54.83 56.603 59.89 56.68 ;
        RECT 54.784 56.649 59.844 56.726 ;
        RECT 54.738 56.695 59.798 56.772 ;
        RECT 54.692 56.741 59.752 56.818 ;
        RECT 54.646 56.787 59.706 56.864 ;
        RECT 54.6 56.833 59.66 56.91 ;
        RECT 54.554 56.879 59.614 56.956 ;
        RECT 54.508 56.925 59.568 57.002 ;
        RECT 54.462 56.971 59.522 57.048 ;
        RECT 54.416 57.017 59.476 57.094 ;
        RECT 54.37 57.063 59.43 57.14 ;
        RECT 54.324 57.109 59.384 57.186 ;
        RECT 54.278 57.155 59.338 57.232 ;
        RECT 54.232 57.201 59.292 57.278 ;
        RECT 54.186 57.247 59.246 57.324 ;
        RECT 54.14 57.293 59.2 57.37 ;
        RECT 54.094 57.339 59.154 57.416 ;
        RECT 54.048 57.385 59.108 57.462 ;
        RECT 54.002 57.431 59.062 57.508 ;
        RECT 53.956 57.477 59.016 57.554 ;
        RECT 53.91 57.523 58.97 57.6 ;
        RECT 53.864 57.569 58.924 57.646 ;
        RECT 53.818 57.615 58.878 57.692 ;
        RECT 53.772 57.661 58.832 57.738 ;
        RECT 53.726 57.707 58.786 57.784 ;
        RECT 53.68 57.753 58.74 57.83 ;
        RECT 53.634 57.799 58.694 57.876 ;
        RECT 53.588 57.845 58.648 57.922 ;
        RECT 53.542 57.891 58.602 57.968 ;
        RECT 53.496 57.937 58.556 58.014 ;
        RECT 53.45 57.983 58.51 58.06 ;
        RECT 53.404 58.029 58.464 58.106 ;
        RECT 53.358 58.075 58.418 58.152 ;
        RECT 53.312 58.121 58.372 58.198 ;
        RECT 53.266 58.167 58.326 58.244 ;
        RECT 53.22 58.213 58.28 58.29 ;
        RECT 53.174 58.259 58.234 58.336 ;
        RECT 53.128 58.305 58.188 58.382 ;
        RECT 53.082 58.351 58.142 58.428 ;
        RECT 53.036 58.397 58.096 58.474 ;
        RECT 52.99 58.443 58.05 58.52 ;
        RECT 52.944 58.489 58.004 58.566 ;
        RECT 52.898 58.535 57.958 58.612 ;
        RECT 52.852 58.581 57.912 58.658 ;
        RECT 52.806 58.627 57.866 58.704 ;
        RECT 52.76 58.673 57.82 58.75 ;
        RECT 52.714 58.719 57.774 58.796 ;
        RECT 52.668 58.765 57.728 58.842 ;
        RECT 52.622 58.811 57.682 58.888 ;
        RECT 52.576 58.857 57.636 58.934 ;
        RECT 52.53 58.903 57.59 58.98 ;
        RECT 52.484 58.949 57.544 59.026 ;
        RECT 52.438 58.995 57.498 59.072 ;
        RECT 52.392 59.041 57.452 59.118 ;
        RECT 52.346 59.087 57.406 59.164 ;
        RECT 52.3 59.133 57.36 59.21 ;
        RECT 52.254 59.179 57.314 59.256 ;
        RECT 52.208 59.225 57.268 59.302 ;
        RECT 52.162 59.271 57.222 59.348 ;
        RECT 52.116 59.317 57.176 59.394 ;
        RECT 52.07 59.363 57.13 59.44 ;
        RECT 52.024 59.409 57.084 59.486 ;
        RECT 51.978 59.455 57.038 59.532 ;
        RECT 51.932 59.501 56.992 59.578 ;
        RECT 51.886 59.547 56.946 59.624 ;
        RECT 51.84 59.593 56.9 59.67 ;
        RECT 51.794 59.639 56.854 59.716 ;
        RECT 51.748 59.685 56.808 59.762 ;
        RECT 51.702 59.731 56.762 59.808 ;
        RECT 51.656 59.777 56.716 59.854 ;
        RECT 51.61 59.823 56.67 59.9 ;
        RECT 51.564 59.869 56.624 59.946 ;
        RECT 51.518 59.915 56.578 59.992 ;
        RECT 51.472 59.961 56.532 60.038 ;
        RECT 51.426 60.007 56.486 60.084 ;
        RECT 51.38 60.053 56.44 60.13 ;
        RECT 51.334 60.099 56.394 60.176 ;
        RECT 51.288 60.145 56.348 60.222 ;
        RECT 51.242 60.191 56.302 60.268 ;
        RECT 51.196 60.237 56.256 60.314 ;
        RECT 51.15 60.283 56.21 60.36 ;
        RECT 51.104 60.329 56.164 60.406 ;
        RECT 51.058 60.375 56.118 60.452 ;
        RECT 51.012 60.421 56.072 60.498 ;
        RECT 50.966 60.467 56.026 60.544 ;
        RECT 50.92 60.513 55.98 60.59 ;
        RECT 50.874 60.559 55.934 60.636 ;
        RECT 50.828 60.605 55.888 60.682 ;
        RECT 50.782 60.651 55.842 60.728 ;
        RECT 50.736 60.697 55.796 60.774 ;
        RECT 50.69 60.743 55.75 60.82 ;
        RECT 50.644 60.789 55.704 60.866 ;
        RECT 50.598 60.835 55.658 60.912 ;
        RECT 50.552 60.881 55.612 60.958 ;
        RECT 50.506 60.927 55.566 61.004 ;
        RECT 50.46 60.973 55.52 61.05 ;
        RECT 50.414 61.019 55.474 61.096 ;
        RECT 50.368 61.065 55.428 61.142 ;
        RECT 50.322 61.111 55.382 61.188 ;
        RECT 50.276 61.157 55.336 61.234 ;
        RECT 50.23 61.203 55.29 61.28 ;
        RECT 50.184 61.249 55.244 61.326 ;
        RECT 50.138 61.295 55.198 61.372 ;
        RECT 50.092 61.341 55.152 61.418 ;
        RECT 50.046 61.387 55.106 61.464 ;
        RECT 50 61.433 55.06 61.51 ;
        RECT 49.954 61.479 55.014 61.556 ;
        RECT 49.908 61.525 54.968 61.602 ;
        RECT 49.862 61.571 54.922 61.648 ;
        RECT 49.816 61.617 54.876 61.694 ;
        RECT 49.77 61.663 54.83 61.74 ;
        RECT 49.724 61.709 54.784 61.786 ;
        RECT 49.678 61.755 54.738 61.832 ;
        RECT 49.632 61.801 54.692 61.878 ;
        RECT 49.586 61.847 54.646 61.924 ;
        RECT 49.54 61.893 54.6 61.97 ;
        RECT 49.494 61.939 54.554 62.016 ;
        RECT 49.448 61.985 54.508 62.062 ;
        RECT 49.402 62.031 54.462 62.108 ;
        RECT 49.356 62.077 54.416 62.154 ;
        RECT 49.31 62.123 54.37 62.2 ;
        RECT 49.264 62.169 54.324 62.246 ;
        RECT 49.218 62.215 54.278 62.292 ;
        RECT 49.172 62.261 54.232 62.338 ;
        RECT 49.126 62.307 54.186 62.384 ;
        RECT 49.08 62.353 54.14 62.43 ;
        RECT 49.034 62.399 54.094 62.476 ;
        RECT 48.988 62.445 54.048 62.522 ;
        RECT 48.942 62.491 54.002 62.568 ;
        RECT 48.85 62.583 53.956 62.614 ;
        RECT 48.896 62.537 53.956 62.614 ;
        RECT 48.838 62.612 53.91 62.66 ;
        RECT 48.792 62.641 53.864 62.706 ;
        RECT 48.746 62.687 53.818 62.752 ;
        RECT 48.7 62.733 53.772 62.798 ;
        RECT 48.654 62.779 53.726 62.844 ;
        RECT 48.608 62.825 53.68 62.89 ;
        RECT 48.562 62.871 53.634 62.936 ;
        RECT 48.516 62.917 53.588 62.982 ;
        RECT 48.47 62.963 53.542 63.028 ;
        RECT 48.424 63.009 53.496 63.074 ;
        RECT 48.378 63.055 53.45 63.12 ;
        RECT 48.332 63.101 53.404 63.166 ;
        RECT 48.286 63.147 53.358 63.212 ;
        RECT 48.24 63.193 53.312 63.258 ;
        RECT 48.194 63.239 53.266 63.304 ;
        RECT 48.148 63.285 53.22 63.35 ;
        RECT 48.102 63.331 53.174 63.396 ;
        RECT 48.056 63.377 53.128 63.442 ;
        RECT 48.01 63.423 53.082 63.488 ;
        RECT 47.964 63.469 53.036 63.534 ;
        RECT 47.918 63.515 52.99 63.58 ;
        RECT 47.872 63.561 52.944 63.626 ;
        RECT 47.826 63.607 52.898 63.672 ;
        RECT 47.78 63.653 52.852 63.718 ;
        RECT 47.734 63.699 52.806 63.764 ;
        RECT 47.688 63.745 52.76 63.81 ;
        RECT 47.642 63.791 52.714 63.856 ;
        RECT 47.596 63.837 52.668 63.902 ;
        RECT 47.55 63.883 52.622 63.948 ;
        RECT 47.504 63.929 52.576 63.994 ;
        RECT 47.458 63.975 52.53 64.04 ;
        RECT 47.412 64.021 52.484 64.086 ;
        RECT 47.366 64.067 52.438 64.132 ;
        RECT 47.32 64.113 52.392 64.178 ;
        RECT 47.274 64.159 52.346 64.224 ;
        RECT 47.228 64.205 52.3 64.27 ;
        RECT 47.182 64.251 52.254 64.316 ;
        RECT 47.136 64.297 52.208 64.362 ;
        RECT 47.09 64.343 52.162 64.408 ;
        RECT 47.044 64.389 52.116 64.454 ;
        RECT 46.998 64.435 52.07 64.5 ;
        RECT 46.952 64.481 52.024 64.546 ;
        RECT 46.906 64.527 51.978 64.592 ;
        RECT 46.86 64.573 51.932 64.638 ;
        RECT 46.814 64.619 51.886 64.684 ;
        RECT 46.768 64.665 51.84 64.73 ;
        RECT 46.722 64.711 51.794 64.776 ;
        RECT 46.676 64.757 51.748 64.822 ;
        RECT 46.63 64.803 51.702 64.868 ;
        RECT 46.584 64.849 51.656 64.914 ;
        RECT 46.538 64.895 51.61 64.96 ;
        RECT 46.492 64.941 51.564 65.006 ;
        RECT 46.446 64.987 51.518 65.052 ;
        RECT 46.4 65.033 51.472 65.098 ;
        RECT 46.354 65.079 51.426 65.144 ;
        RECT 46.308 65.125 51.38 65.19 ;
        RECT 46.262 65.171 51.334 65.236 ;
        RECT 46.216 65.217 51.288 65.282 ;
        RECT 46.17 65.263 51.242 65.328 ;
        RECT 46.124 65.309 51.196 65.374 ;
        RECT 46.078 65.355 51.15 65.42 ;
        RECT 46.032 65.401 51.104 65.466 ;
        RECT 45.986 65.447 51.058 65.512 ;
        RECT 45.94 65.493 51.012 65.558 ;
        RECT 45.894 65.539 50.966 65.604 ;
        RECT 45.848 65.585 50.92 65.65 ;
        RECT 45.802 65.631 50.874 65.696 ;
        RECT 45.756 65.677 50.828 65.742 ;
        RECT 45.71 65.723 50.782 65.788 ;
        RECT 45.664 65.769 50.736 65.834 ;
        RECT 45.618 65.815 50.69 65.88 ;
        RECT 45.572 65.861 50.644 65.926 ;
        RECT 45.526 65.907 50.598 65.972 ;
        RECT 45.48 65.953 50.552 66.018 ;
        RECT 45.434 65.999 50.506 66.064 ;
        RECT 45.388 66.045 50.46 66.11 ;
        RECT 45.342 66.091 50.414 66.156 ;
        RECT 45.296 66.137 50.368 66.202 ;
        RECT 45.25 66.183 50.322 66.248 ;
        RECT 45.25 66.183 50.276 66.294 ;
        RECT 45.25 66.183 50.23 66.34 ;
        RECT 45.25 66.183 50.184 66.386 ;
        RECT 45.25 66.183 50.138 66.432 ;
        RECT 45.25 66.183 50.092 66.478 ;
        RECT 45.25 66.183 50.046 66.524 ;
        RECT 45.25 66.183 50 66.57 ;
        RECT 45.25 66.183 49.954 66.616 ;
        RECT 45.25 66.183 49.908 66.662 ;
        RECT 45.25 66.183 49.862 66.708 ;
        RECT 45.25 66.183 49.816 66.754 ;
        RECT 45.25 66.183 49.77 66.8 ;
        RECT 45.25 66.183 49.724 66.846 ;
        RECT 45.25 66.183 49.678 66.892 ;
        RECT 45.25 66.183 49.632 66.938 ;
        RECT 45.25 66.183 49.586 66.984 ;
        RECT 45.25 66.183 49.54 67.03 ;
        RECT 45.25 66.183 49.494 67.076 ;
        RECT 45.25 66.183 49.448 67.122 ;
        RECT 45.25 66.183 49.402 67.168 ;
        RECT 45.25 66.183 49.356 67.214 ;
        RECT 45.25 66.183 49.31 67.26 ;
        RECT 45.25 66.183 49.264 67.306 ;
        RECT 45.25 66.183 49.218 67.352 ;
        RECT 45.25 66.183 49.172 67.398 ;
        RECT 45.25 66.183 49.126 67.444 ;
        RECT 45.25 66.183 49.08 67.49 ;
        RECT 45.25 66.183 49.034 67.536 ;
        RECT 45.25 66.183 48.988 67.582 ;
        RECT 45.25 66.183 48.942 67.628 ;
        RECT 45.25 66.183 48.896 67.674 ;
        RECT 45.25 66.183 48.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 62.504 42.281 62.55 47.372 ;
        RECT 57.444 47.341 62.504 47.418 ;
        RECT 61.032 43.753 80 44.15 ;
        RECT 62.458 42.327 62.504 47.418 ;
        RECT 57.398 47.387 62.458 47.464 ;
        RECT 61.078 43.707 80 44.15 ;
        RECT 62.412 42.373 62.458 47.464 ;
        RECT 57.352 47.433 62.412 47.51 ;
        RECT 61.124 43.661 80 44.15 ;
        RECT 62.366 42.419 62.412 47.51 ;
        RECT 57.306 47.479 62.366 47.556 ;
        RECT 61.17 43.615 80 44.15 ;
        RECT 62.32 42.465 62.366 47.556 ;
        RECT 57.26 47.525 62.32 47.602 ;
        RECT 61.216 43.569 80 44.15 ;
        RECT 62.274 42.511 62.32 47.602 ;
        RECT 57.214 47.571 62.274 47.648 ;
        RECT 61.262 43.523 80 44.15 ;
        RECT 62.228 42.557 62.274 47.648 ;
        RECT 57.168 47.617 62.228 47.694 ;
        RECT 61.308 43.477 80 44.15 ;
        RECT 62.182 42.603 62.228 47.694 ;
        RECT 57.122 47.663 62.182 47.74 ;
        RECT 61.354 43.431 80 44.15 ;
        RECT 62.136 42.649 62.182 47.74 ;
        RECT 57.076 47.709 62.136 47.786 ;
        RECT 61.4 43.385 80 44.15 ;
        RECT 62.09 42.695 62.136 47.786 ;
        RECT 57.03 47.755 62.09 47.832 ;
        RECT 61.446 43.339 80 44.15 ;
        RECT 62.044 42.741 62.09 47.832 ;
        RECT 56.984 47.801 62.044 47.878 ;
        RECT 61.492 43.293 80 44.15 ;
        RECT 61.998 42.787 62.044 47.878 ;
        RECT 56.938 47.847 61.998 47.924 ;
        RECT 61.538 43.247 80 44.15 ;
        RECT 61.952 42.833 61.998 47.924 ;
        RECT 56.892 47.893 61.952 47.97 ;
        RECT 61.584 43.201 80 44.15 ;
        RECT 61.906 42.879 61.952 47.97 ;
        RECT 56.846 47.939 61.906 48.016 ;
        RECT 61.63 43.155 80 44.15 ;
        RECT 61.86 42.925 61.906 48.016 ;
        RECT 56.8 47.985 61.86 48.062 ;
        RECT 61.676 43.109 80 44.15 ;
        RECT 61.814 42.971 61.86 48.062 ;
        RECT 56.754 48.031 61.814 48.108 ;
        RECT 61.722 43.063 80 44.15 ;
        RECT 61.768 43.017 61.814 48.108 ;
        RECT 56.708 48.077 61.768 48.154 ;
        RECT 56.662 48.123 61.722 48.2 ;
        RECT 56.616 48.169 61.676 48.246 ;
        RECT 56.57 48.215 61.63 48.292 ;
        RECT 56.524 48.261 61.584 48.338 ;
        RECT 56.478 48.307 61.538 48.384 ;
        RECT 56.432 48.353 61.492 48.43 ;
        RECT 56.386 48.399 61.446 48.476 ;
        RECT 56.34 48.445 61.4 48.522 ;
        RECT 56.294 48.491 61.354 48.568 ;
        RECT 56.248 48.537 61.308 48.614 ;
        RECT 56.202 48.583 61.262 48.66 ;
        RECT 56.156 48.629 61.216 48.706 ;
        RECT 56.11 48.675 61.17 48.752 ;
        RECT 56.064 48.721 61.124 48.798 ;
        RECT 56.018 48.767 61.078 48.844 ;
        RECT 55.972 48.813 61.032 48.89 ;
        RECT 55.926 48.859 60.986 48.936 ;
        RECT 55.88 48.905 60.94 48.982 ;
        RECT 55.834 48.951 60.894 49.028 ;
        RECT 55.788 48.997 60.848 49.074 ;
        RECT 55.742 49.043 60.802 49.12 ;
        RECT 55.696 49.089 60.756 49.166 ;
        RECT 55.65 49.135 60.71 49.212 ;
        RECT 55.604 49.181 60.664 49.258 ;
        RECT 55.558 49.227 60.618 49.304 ;
        RECT 55.512 49.273 60.572 49.35 ;
        RECT 55.466 49.319 60.526 49.396 ;
        RECT 55.42 49.365 60.48 49.442 ;
        RECT 55.374 49.411 60.434 49.488 ;
        RECT 55.328 49.457 60.388 49.534 ;
        RECT 55.282 49.503 60.342 49.58 ;
        RECT 55.236 49.549 60.296 49.626 ;
        RECT 55.19 49.595 60.25 49.672 ;
        RECT 55.144 49.641 60.204 49.718 ;
        RECT 55.098 49.687 60.158 49.764 ;
        RECT 55.052 49.733 60.112 49.81 ;
        RECT 55.006 49.779 60.066 49.856 ;
        RECT 54.96 49.825 60.02 49.902 ;
        RECT 54.914 49.871 59.974 49.948 ;
        RECT 54.868 49.917 59.928 49.994 ;
        RECT 54.822 49.963 59.882 50.04 ;
        RECT 54.776 50.009 59.836 50.086 ;
        RECT 54.73 50.055 59.79 50.132 ;
        RECT 54.684 50.101 59.744 50.178 ;
        RECT 54.638 50.147 59.698 50.224 ;
        RECT 54.592 50.193 59.652 50.27 ;
        RECT 54.546 50.239 59.606 50.316 ;
        RECT 54.5 50.285 59.56 50.362 ;
        RECT 54.454 50.331 59.514 50.408 ;
        RECT 54.408 50.377 59.468 50.454 ;
        RECT 54.362 50.423 59.422 50.5 ;
        RECT 54.316 50.469 59.376 50.546 ;
        RECT 54.27 50.515 59.33 50.592 ;
        RECT 54.224 50.561 59.284 50.638 ;
        RECT 54.178 50.607 59.238 50.684 ;
        RECT 54.132 50.653 59.192 50.73 ;
        RECT 54.086 50.699 59.146 50.776 ;
        RECT 54.04 50.745 59.1 50.822 ;
        RECT 53.994 50.791 59.054 50.868 ;
        RECT 53.948 50.837 59.008 50.914 ;
        RECT 53.902 50.883 58.962 50.96 ;
        RECT 53.856 50.929 58.916 51.006 ;
        RECT 53.81 50.975 58.87 51.052 ;
        RECT 53.764 51.021 58.824 51.098 ;
        RECT 53.718 51.067 58.778 51.144 ;
        RECT 53.672 51.113 58.732 51.19 ;
        RECT 53.626 51.159 58.686 51.236 ;
        RECT 53.58 51.205 58.64 51.282 ;
        RECT 53.534 51.251 58.594 51.328 ;
        RECT 53.488 51.297 58.548 51.374 ;
        RECT 53.442 51.343 58.502 51.42 ;
        RECT 53.396 51.389 58.456 51.466 ;
        RECT 53.35 51.435 58.41 51.512 ;
        RECT 53.304 51.481 58.364 51.558 ;
        RECT 53.258 51.527 58.318 51.604 ;
        RECT 53.212 51.573 58.272 51.65 ;
        RECT 53.166 51.619 58.226 51.696 ;
        RECT 53.12 51.665 58.18 51.742 ;
        RECT 53.074 51.711 58.134 51.788 ;
        RECT 53.028 51.757 58.088 51.834 ;
        RECT 52.982 51.803 58.042 51.88 ;
        RECT 52.936 51.849 57.996 51.926 ;
        RECT 52.89 51.895 57.95 51.972 ;
        RECT 52.844 51.941 57.904 52.018 ;
        RECT 52.798 51.987 57.858 52.064 ;
        RECT 52.752 52.033 57.812 52.11 ;
        RECT 52.706 52.079 57.766 52.156 ;
        RECT 52.66 52.125 57.72 52.202 ;
        RECT 52.614 52.171 57.674 52.248 ;
        RECT 52.568 52.217 57.628 52.294 ;
        RECT 52.522 52.263 57.582 52.34 ;
        RECT 52.476 52.309 57.536 52.386 ;
        RECT 52.43 52.355 57.49 52.432 ;
        RECT 52.384 52.401 57.444 52.478 ;
        RECT 52.338 52.447 57.398 52.524 ;
        RECT 52.292 52.493 57.352 52.57 ;
        RECT 52.246 52.539 57.306 52.616 ;
        RECT 52.2 52.585 57.26 52.662 ;
        RECT 52.154 52.631 57.214 52.708 ;
        RECT 52.108 52.677 57.168 52.754 ;
        RECT 52.062 52.723 57.122 52.8 ;
        RECT 52.016 52.769 57.076 52.846 ;
        RECT 51.97 52.815 57.03 52.892 ;
        RECT 51.924 52.861 56.984 52.938 ;
        RECT 51.878 52.907 56.938 52.984 ;
        RECT 51.832 52.953 56.892 53.03 ;
        RECT 51.786 52.999 56.846 53.076 ;
        RECT 51.74 53.045 56.8 53.122 ;
        RECT 51.694 53.091 56.754 53.168 ;
        RECT 51.648 53.137 56.708 53.214 ;
        RECT 51.602 53.183 56.662 53.26 ;
        RECT 51.556 53.229 56.616 53.306 ;
        RECT 51.51 53.275 56.57 53.352 ;
        RECT 51.464 53.321 56.524 53.398 ;
        RECT 51.418 53.367 56.478 53.444 ;
        RECT 51.372 53.413 56.432 53.49 ;
        RECT 51.326 53.459 56.386 53.536 ;
        RECT 51.28 53.505 56.34 53.582 ;
        RECT 51.234 53.551 56.294 53.628 ;
        RECT 51.188 53.597 56.248 53.674 ;
        RECT 51.142 53.643 56.202 53.72 ;
        RECT 51.096 53.689 56.156 53.766 ;
        RECT 51.05 53.735 56.11 53.812 ;
        RECT 51.004 53.781 56.064 53.858 ;
        RECT 50.958 53.827 56.018 53.904 ;
        RECT 50.912 53.873 55.972 53.95 ;
        RECT 50.866 53.919 55.926 53.996 ;
        RECT 50.82 53.965 55.88 54.042 ;
        RECT 50.774 54.011 55.834 54.088 ;
        RECT 50.728 54.057 55.788 54.134 ;
        RECT 50.682 54.103 55.742 54.18 ;
        RECT 50.636 54.149 55.696 54.226 ;
        RECT 50.59 54.195 55.65 54.272 ;
        RECT 50.544 54.241 55.604 54.318 ;
        RECT 50.498 54.287 55.558 54.364 ;
        RECT 50.452 54.333 55.512 54.41 ;
        RECT 50.406 54.379 55.466 54.456 ;
        RECT 50.36 54.425 55.42 54.502 ;
        RECT 50.314 54.471 55.374 54.548 ;
        RECT 50.268 54.517 55.328 54.594 ;
        RECT 50.222 54.563 55.282 54.64 ;
        RECT 50.176 54.609 55.236 54.686 ;
        RECT 50.13 54.655 55.19 54.732 ;
        RECT 50.084 54.701 55.144 54.778 ;
        RECT 50.038 54.747 55.098 54.824 ;
        RECT 49.992 54.793 55.052 54.87 ;
        RECT 49.946 54.839 55.006 54.916 ;
        RECT 49.9 54.885 54.96 54.962 ;
        RECT 49.854 54.931 54.914 55.008 ;
        RECT 49.808 54.977 54.868 55.054 ;
        RECT 49.762 55.023 54.822 55.1 ;
        RECT 49.716 55.069 54.776 55.146 ;
        RECT 49.67 55.115 54.73 55.192 ;
        RECT 49.624 55.161 54.684 55.238 ;
        RECT 49.578 55.207 54.638 55.284 ;
        RECT 49.532 55.253 54.592 55.33 ;
        RECT 49.486 55.299 54.546 55.376 ;
        RECT 49.44 55.345 54.5 55.422 ;
        RECT 49.394 55.391 54.454 55.468 ;
        RECT 49.348 55.437 54.408 55.514 ;
        RECT 49.302 55.483 54.362 55.56 ;
        RECT 49.256 55.529 54.316 55.606 ;
        RECT 49.21 55.575 54.27 55.652 ;
        RECT 49.164 55.621 54.224 55.698 ;
        RECT 49.118 55.667 54.178 55.744 ;
        RECT 49.072 55.713 54.132 55.79 ;
        RECT 49.026 55.759 54.086 55.836 ;
        RECT 48.98 55.805 54.04 55.882 ;
        RECT 48.934 55.851 53.994 55.928 ;
        RECT 48.888 55.897 53.948 55.974 ;
        RECT 48.842 55.943 53.902 56.02 ;
        RECT 48.796 55.989 53.856 56.066 ;
        RECT 48.75 56.035 53.81 56.112 ;
        RECT 48.704 56.081 53.764 56.158 ;
        RECT 48.658 56.127 53.718 56.204 ;
        RECT 48.612 56.173 53.672 56.25 ;
        RECT 48.566 56.219 53.626 56.296 ;
        RECT 48.52 56.265 53.58 56.342 ;
        RECT 48.474 56.311 53.534 56.388 ;
        RECT 48.428 56.357 53.488 56.434 ;
        RECT 48.382 56.403 53.442 56.48 ;
        RECT 48.336 56.449 53.396 56.526 ;
        RECT 48.29 56.495 53.35 56.572 ;
        RECT 48.244 56.541 53.304 56.618 ;
        RECT 48.198 56.587 53.258 56.664 ;
        RECT 48.152 56.633 53.212 56.71 ;
        RECT 48.106 56.679 53.166 56.756 ;
        RECT 48.06 56.725 53.12 56.802 ;
        RECT 48.014 56.771 53.074 56.848 ;
        RECT 47.968 56.817 53.028 56.894 ;
        RECT 47.922 56.863 52.982 56.94 ;
        RECT 47.876 56.909 52.936 56.986 ;
        RECT 47.83 56.955 52.89 57.032 ;
        RECT 47.784 57.001 52.844 57.078 ;
        RECT 47.738 57.047 52.798 57.124 ;
        RECT 47.692 57.093 52.752 57.17 ;
        RECT 47.646 57.139 52.706 57.216 ;
        RECT 47.6 57.185 52.66 57.262 ;
        RECT 47.554 57.231 52.614 57.308 ;
        RECT 47.508 57.277 52.568 57.354 ;
        RECT 47.462 57.323 52.522 57.4 ;
        RECT 47.416 57.369 52.476 57.446 ;
        RECT 47.37 57.415 52.43 57.492 ;
        RECT 47.324 57.461 52.384 57.538 ;
        RECT 47.278 57.507 52.338 57.584 ;
        RECT 47.232 57.553 52.292 57.63 ;
        RECT 47.186 57.599 52.246 57.676 ;
        RECT 47.14 57.645 52.2 57.722 ;
        RECT 47.094 57.691 52.154 57.768 ;
        RECT 47.048 57.737 52.108 57.814 ;
        RECT 47.002 57.783 52.062 57.86 ;
        RECT 46.956 57.829 52.016 57.906 ;
        RECT 46.91 57.875 51.97 57.952 ;
        RECT 46.864 57.921 51.924 57.998 ;
        RECT 46.818 57.967 51.878 58.044 ;
        RECT 46.772 58.013 51.832 58.09 ;
        RECT 46.726 58.059 51.786 58.136 ;
        RECT 46.68 58.105 51.74 58.182 ;
        RECT 46.634 58.151 51.694 58.228 ;
        RECT 46.588 58.197 51.648 58.274 ;
        RECT 46.542 58.243 51.602 58.32 ;
        RECT 46.496 58.289 51.556 58.366 ;
        RECT 46.45 58.335 51.51 58.412 ;
        RECT 46.404 58.381 51.464 58.458 ;
        RECT 46.358 58.427 51.418 58.504 ;
        RECT 46.312 58.473 51.372 58.55 ;
        RECT 46.266 58.519 51.326 58.596 ;
        RECT 46.22 58.565 51.28 58.642 ;
        RECT 46.174 58.611 51.234 58.688 ;
        RECT 46.128 58.657 51.188 58.734 ;
        RECT 46.082 58.703 51.142 58.78 ;
        RECT 46.036 58.749 51.096 58.826 ;
        RECT 45.99 58.795 51.05 58.872 ;
        RECT 45.944 58.841 51.004 58.918 ;
        RECT 45.898 58.887 50.958 58.964 ;
        RECT 45.852 58.933 50.912 59.01 ;
        RECT 45.806 58.979 50.866 59.056 ;
        RECT 45.76 59.025 50.82 59.102 ;
        RECT 45.714 59.071 50.774 59.148 ;
        RECT 45.668 59.117 50.728 59.194 ;
        RECT 45.622 59.163 50.682 59.24 ;
        RECT 45.576 59.209 50.636 59.286 ;
        RECT 45.53 59.255 50.59 59.332 ;
        RECT 45.484 59.301 50.544 59.378 ;
        RECT 45.438 59.347 50.498 59.424 ;
        RECT 45.392 59.393 50.452 59.47 ;
        RECT 45.346 59.439 50.406 59.516 ;
        RECT 45.3 59.485 50.36 59.562 ;
        RECT 45.254 59.531 50.314 59.608 ;
        RECT 45.208 59.577 50.268 59.654 ;
        RECT 45.162 59.623 50.222 59.7 ;
        RECT 45.116 59.669 50.176 59.746 ;
        RECT 45.07 59.715 50.13 59.792 ;
        RECT 45.024 59.761 50.084 59.838 ;
        RECT 44.978 59.807 50.038 59.884 ;
        RECT 44.932 59.853 49.992 59.93 ;
        RECT 44.886 59.899 49.946 59.976 ;
        RECT 44.84 59.945 49.9 60.022 ;
        RECT 44.794 59.991 49.854 60.068 ;
        RECT 44.748 60.037 49.808 60.114 ;
        RECT 44.702 60.083 49.762 60.16 ;
        RECT 44.656 60.129 49.716 60.206 ;
        RECT 44.61 60.175 49.67 60.252 ;
        RECT 44.564 60.221 49.624 60.298 ;
        RECT 44.518 60.267 49.578 60.344 ;
        RECT 44.472 60.313 49.532 60.39 ;
        RECT 44.426 60.359 49.486 60.436 ;
        RECT 44.38 60.405 49.44 60.482 ;
        RECT 44.334 60.451 49.394 60.528 ;
        RECT 44.288 60.497 49.348 60.574 ;
        RECT 44.242 60.543 49.302 60.62 ;
        RECT 44.15 60.635 49.256 60.666 ;
        RECT 44.196 60.589 49.256 60.666 ;
        RECT 44.138 60.664 49.21 60.712 ;
        RECT 44.092 60.693 49.164 60.758 ;
        RECT 44.046 60.739 49.118 60.804 ;
        RECT 44 60.785 49.072 60.85 ;
        RECT 43.954 60.831 49.026 60.896 ;
        RECT 43.908 60.877 48.98 60.942 ;
        RECT 43.862 60.923 48.934 60.988 ;
        RECT 43.816 60.969 48.888 61.034 ;
        RECT 43.77 61.015 48.842 61.08 ;
        RECT 43.724 61.061 48.796 61.126 ;
        RECT 43.678 61.107 48.75 61.172 ;
        RECT 43.632 61.153 48.704 61.218 ;
        RECT 43.586 61.199 48.658 61.264 ;
        RECT 43.54 61.245 48.612 61.31 ;
        RECT 43.494 61.291 48.566 61.356 ;
        RECT 43.448 61.337 48.52 61.402 ;
        RECT 43.402 61.383 48.474 61.448 ;
        RECT 43.356 61.429 48.428 61.494 ;
        RECT 43.31 61.475 48.382 61.54 ;
        RECT 43.264 61.521 48.336 61.586 ;
        RECT 43.218 61.567 48.29 61.632 ;
        RECT 43.172 61.613 48.244 61.678 ;
        RECT 43.126 61.659 48.198 61.724 ;
        RECT 43.08 61.705 48.152 61.77 ;
        RECT 43.034 61.751 48.106 61.816 ;
        RECT 42.988 61.797 48.06 61.862 ;
        RECT 42.942 61.843 48.014 61.908 ;
        RECT 42.896 61.889 47.968 61.954 ;
        RECT 42.85 61.935 47.922 62 ;
        RECT 42.804 61.981 47.876 62.046 ;
        RECT 42.758 62.027 47.83 62.092 ;
        RECT 42.712 62.073 47.784 62.138 ;
        RECT 42.666 62.119 47.738 62.184 ;
        RECT 42.62 62.165 47.692 62.23 ;
        RECT 42.574 62.211 47.646 62.276 ;
        RECT 42.528 62.257 47.6 62.322 ;
        RECT 42.482 62.303 47.554 62.368 ;
        RECT 42.436 62.349 47.508 62.414 ;
        RECT 42.39 62.395 47.462 62.46 ;
        RECT 42.344 62.441 47.416 62.506 ;
        RECT 42.298 62.487 47.37 62.552 ;
        RECT 42.252 62.533 47.324 62.598 ;
        RECT 42.206 62.579 47.278 62.644 ;
        RECT 42.16 62.625 47.232 62.69 ;
        RECT 42.114 62.671 47.186 62.736 ;
        RECT 42.068 62.717 47.14 62.782 ;
        RECT 42.022 62.763 47.094 62.828 ;
        RECT 41.976 62.809 47.048 62.874 ;
        RECT 41.93 62.855 47.002 62.92 ;
        RECT 41.884 62.901 46.956 62.966 ;
        RECT 41.838 62.947 46.91 63.012 ;
        RECT 41.792 62.993 46.864 63.058 ;
        RECT 41.746 63.039 46.818 63.104 ;
        RECT 41.7 63.085 46.772 63.15 ;
        RECT 41.654 63.131 46.726 63.196 ;
        RECT 41.608 63.177 46.68 63.242 ;
        RECT 41.562 63.223 46.634 63.288 ;
        RECT 41.516 63.269 46.588 63.334 ;
        RECT 41.47 63.315 46.542 63.38 ;
        RECT 41.424 63.361 46.496 63.426 ;
        RECT 41.378 63.407 46.45 63.472 ;
        RECT 41.332 63.453 46.404 63.518 ;
        RECT 41.286 63.499 46.358 63.564 ;
        RECT 41.24 63.545 46.312 63.61 ;
        RECT 41.194 63.591 46.266 63.656 ;
        RECT 41.148 63.637 46.22 63.702 ;
        RECT 41.102 63.683 46.174 63.748 ;
        RECT 41.056 63.729 46.128 63.794 ;
        RECT 41.01 63.775 46.082 63.84 ;
        RECT 40.964 63.821 46.036 63.886 ;
        RECT 40.918 63.867 45.99 63.932 ;
        RECT 40.872 63.913 45.944 63.978 ;
        RECT 40.826 63.959 45.898 64.024 ;
        RECT 40.78 64.005 45.852 64.07 ;
        RECT 40.734 64.051 45.806 64.116 ;
        RECT 40.688 64.097 45.76 64.162 ;
        RECT 40.642 64.143 45.714 64.208 ;
        RECT 40.596 64.189 45.668 64.254 ;
        RECT 40.55 64.235 45.622 64.3 ;
        RECT 40.55 64.235 45.576 64.346 ;
        RECT 40.55 64.235 45.53 64.392 ;
        RECT 40.55 64.235 45.484 64.438 ;
        RECT 40.55 64.235 45.438 64.484 ;
        RECT 40.55 64.235 45.392 64.53 ;
        RECT 40.55 64.235 45.346 64.576 ;
        RECT 40.55 64.235 45.3 64.622 ;
        RECT 40.55 64.235 45.254 64.668 ;
        RECT 40.55 64.235 45.208 64.714 ;
        RECT 40.55 64.235 45.162 64.76 ;
        RECT 40.55 64.235 45.116 64.806 ;
        RECT 40.55 64.235 45.07 64.852 ;
        RECT 40.55 64.235 45.024 64.898 ;
        RECT 40.55 64.235 44.978 64.944 ;
        RECT 40.55 64.235 44.932 64.99 ;
        RECT 40.55 64.235 44.886 65.036 ;
        RECT 40.55 64.235 44.84 65.082 ;
        RECT 40.55 64.235 44.794 65.128 ;
        RECT 40.55 64.235 44.748 65.174 ;
        RECT 40.55 64.235 44.702 65.22 ;
        RECT 40.55 64.235 44.656 65.266 ;
        RECT 40.55 64.235 44.61 65.312 ;
        RECT 40.55 64.235 44.564 65.358 ;
        RECT 40.55 64.235 44.518 65.404 ;
        RECT 40.55 64.235 44.472 65.45 ;
        RECT 40.55 64.235 44.426 65.496 ;
        RECT 40.55 64.235 44.38 65.542 ;
        RECT 40.55 64.235 44.334 65.588 ;
        RECT 40.55 64.235 44.288 65.634 ;
        RECT 40.55 64.235 44.242 65.68 ;
        RECT 40.55 64.235 44.196 65.726 ;
        RECT 40.55 64.235 44.15 80 ;
        RECT 64.258 40.55 80 44.15 ;
        RECT 60.664 44.121 65.749 44.16 ;
        RECT 59.192 45.593 64.258 45.644 ;
        RECT 59.238 45.547 64.304 45.618 ;
        RECT 64.252 40.553 64.258 45.644 ;
        RECT 59.284 45.501 64.35 45.572 ;
        RECT 64.206 40.579 64.252 45.67 ;
        RECT 59.146 45.639 64.206 45.716 ;
        RECT 59.33 45.455 64.396 45.526 ;
        RECT 64.16 40.625 64.206 45.716 ;
        RECT 59.1 45.685 64.16 45.762 ;
        RECT 59.376 45.409 64.442 45.48 ;
        RECT 64.114 40.671 64.16 45.762 ;
        RECT 59.054 45.731 64.114 45.808 ;
        RECT 59.422 45.363 64.488 45.434 ;
        RECT 64.068 40.717 64.114 45.808 ;
        RECT 59.008 45.777 64.068 45.854 ;
        RECT 59.468 45.317 64.534 45.388 ;
        RECT 64.022 40.763 64.068 45.854 ;
        RECT 58.962 45.823 64.022 45.9 ;
        RECT 59.514 45.271 64.58 45.342 ;
        RECT 63.976 40.809 64.022 45.9 ;
        RECT 58.916 45.869 63.976 45.946 ;
        RECT 59.56 45.225 64.626 45.296 ;
        RECT 63.93 40.855 63.976 45.946 ;
        RECT 58.87 45.915 63.93 45.992 ;
        RECT 59.606 45.179 64.672 45.25 ;
        RECT 63.884 40.901 63.93 45.992 ;
        RECT 58.824 45.961 63.884 46.038 ;
        RECT 59.652 45.133 64.718 45.204 ;
        RECT 63.838 40.947 63.884 46.038 ;
        RECT 58.778 46.007 63.838 46.084 ;
        RECT 59.698 45.087 64.764 45.158 ;
        RECT 63.792 40.993 63.838 46.084 ;
        RECT 58.732 46.053 63.792 46.13 ;
        RECT 59.744 45.041 64.81 45.112 ;
        RECT 63.746 41.039 63.792 46.13 ;
        RECT 58.686 46.099 63.746 46.176 ;
        RECT 59.79 44.995 64.856 45.066 ;
        RECT 63.7 41.085 63.746 46.176 ;
        RECT 58.64 46.145 63.7 46.222 ;
        RECT 59.836 44.949 64.902 45.02 ;
        RECT 63.654 41.131 63.7 46.222 ;
        RECT 58.594 46.191 63.654 46.268 ;
        RECT 59.882 44.903 64.948 44.974 ;
        RECT 63.608 41.177 63.654 46.268 ;
        RECT 58.548 46.237 63.608 46.314 ;
        RECT 59.928 44.857 64.994 44.928 ;
        RECT 63.562 41.223 63.608 46.314 ;
        RECT 58.502 46.283 63.562 46.36 ;
        RECT 59.974 44.811 65.04 44.882 ;
        RECT 63.516 41.269 63.562 46.36 ;
        RECT 58.456 46.329 63.516 46.406 ;
        RECT 60.02 44.765 65.086 44.836 ;
        RECT 63.47 41.315 63.516 46.406 ;
        RECT 58.41 46.375 63.47 46.452 ;
        RECT 60.066 44.719 65.132 44.79 ;
        RECT 63.424 41.361 63.47 46.452 ;
        RECT 58.364 46.421 63.424 46.498 ;
        RECT 60.112 44.673 65.178 44.744 ;
        RECT 63.378 41.407 63.424 46.498 ;
        RECT 58.318 46.467 63.378 46.544 ;
        RECT 60.158 44.627 65.224 44.698 ;
        RECT 63.332 41.453 63.378 46.544 ;
        RECT 58.272 46.513 63.332 46.59 ;
        RECT 60.204 44.581 65.27 44.652 ;
        RECT 63.286 41.499 63.332 46.59 ;
        RECT 58.226 46.559 63.286 46.636 ;
        RECT 60.25 44.535 65.316 44.606 ;
        RECT 63.24 41.545 63.286 46.636 ;
        RECT 58.18 46.605 63.24 46.682 ;
        RECT 60.296 44.489 65.362 44.56 ;
        RECT 63.194 41.591 63.24 46.682 ;
        RECT 58.134 46.651 63.194 46.728 ;
        RECT 60.342 44.443 65.408 44.514 ;
        RECT 63.148 41.637 63.194 46.728 ;
        RECT 58.088 46.697 63.148 46.774 ;
        RECT 60.388 44.397 65.454 44.468 ;
        RECT 63.102 41.683 63.148 46.774 ;
        RECT 58.042 46.743 63.102 46.82 ;
        RECT 60.434 44.351 65.5 44.422 ;
        RECT 63.056 41.729 63.102 46.82 ;
        RECT 57.996 46.789 63.056 46.866 ;
        RECT 60.48 44.305 65.546 44.376 ;
        RECT 63.01 41.775 63.056 46.866 ;
        RECT 57.95 46.835 63.01 46.912 ;
        RECT 60.526 44.259 65.592 44.33 ;
        RECT 62.964 41.821 63.01 46.912 ;
        RECT 57.904 46.881 62.964 46.958 ;
        RECT 60.572 44.213 65.638 44.284 ;
        RECT 62.918 41.867 62.964 46.958 ;
        RECT 57.858 46.927 62.918 47.004 ;
        RECT 60.618 44.167 65.684 44.238 ;
        RECT 62.872 41.913 62.918 47.004 ;
        RECT 57.812 46.973 62.872 47.05 ;
        RECT 60.664 44.121 65.73 44.192 ;
        RECT 62.826 41.959 62.872 47.05 ;
        RECT 57.766 47.019 62.826 47.096 ;
        RECT 60.71 44.075 80 44.15 ;
        RECT 62.78 42.005 62.826 47.096 ;
        RECT 57.72 47.065 62.78 47.142 ;
        RECT 60.756 44.029 80 44.15 ;
        RECT 62.734 42.051 62.78 47.142 ;
        RECT 57.674 47.111 62.734 47.188 ;
        RECT 60.802 43.983 80 44.15 ;
        RECT 62.688 42.097 62.734 47.188 ;
        RECT 57.628 47.157 62.688 47.234 ;
        RECT 60.848 43.937 80 44.15 ;
        RECT 62.642 42.143 62.688 47.234 ;
        RECT 57.582 47.203 62.642 47.28 ;
        RECT 60.894 43.891 80 44.15 ;
        RECT 62.596 42.189 62.642 47.28 ;
        RECT 57.536 47.249 62.596 47.326 ;
        RECT 60.94 43.845 80 44.15 ;
        RECT 62.55 42.235 62.596 47.326 ;
        RECT 57.49 47.295 62.55 47.372 ;
        RECT 60.986 43.799 80 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 68.968 55.761 69.014 60.852 ;
        RECT 63.908 60.821 68.968 60.898 ;
        RECT 66.208 58.521 71.298 58.568 ;
        RECT 68.922 55.807 68.968 60.898 ;
        RECT 63.862 60.867 68.922 60.944 ;
        RECT 66.254 58.475 71.344 58.522 ;
        RECT 68.876 55.853 68.922 60.944 ;
        RECT 63.816 60.913 68.876 60.99 ;
        RECT 66.3 58.429 71.39 58.476 ;
        RECT 68.83 55.899 68.876 60.99 ;
        RECT 63.77 60.959 68.83 61.036 ;
        RECT 66.346 58.383 71.436 58.43 ;
        RECT 68.784 55.945 68.83 61.036 ;
        RECT 63.724 61.005 68.784 61.082 ;
        RECT 66.392 58.337 71.482 58.384 ;
        RECT 68.738 55.991 68.784 61.082 ;
        RECT 63.678 61.051 68.738 61.128 ;
        RECT 66.438 58.291 71.528 58.338 ;
        RECT 68.692 56.037 68.738 61.128 ;
        RECT 63.632 61.097 68.692 61.174 ;
        RECT 66.484 58.245 71.574 58.292 ;
        RECT 68.646 56.083 68.692 61.174 ;
        RECT 63.586 61.143 68.646 61.22 ;
        RECT 66.53 58.199 80 58.25 ;
        RECT 68.6 56.129 68.646 61.22 ;
        RECT 63.54 61.189 68.6 61.266 ;
        RECT 66.576 58.153 80 58.25 ;
        RECT 68.554 56.175 68.6 61.266 ;
        RECT 63.494 61.235 68.554 61.312 ;
        RECT 66.622 58.107 80 58.25 ;
        RECT 68.508 56.221 68.554 61.312 ;
        RECT 63.448 61.281 68.508 61.358 ;
        RECT 66.668 58.061 80 58.25 ;
        RECT 68.462 56.267 68.508 61.358 ;
        RECT 63.402 61.327 68.462 61.404 ;
        RECT 66.714 58.015 80 58.25 ;
        RECT 68.416 56.313 68.462 61.404 ;
        RECT 63.356 61.373 68.416 61.45 ;
        RECT 66.76 57.969 80 58.25 ;
        RECT 68.37 56.359 68.416 61.45 ;
        RECT 63.31 61.419 68.37 61.496 ;
        RECT 66.806 57.923 80 58.25 ;
        RECT 68.324 56.405 68.37 61.496 ;
        RECT 63.264 61.465 68.324 61.542 ;
        RECT 66.852 57.877 80 58.25 ;
        RECT 68.278 56.451 68.324 61.542 ;
        RECT 63.218 61.511 68.278 61.588 ;
        RECT 66.898 57.831 80 58.25 ;
        RECT 68.232 56.497 68.278 61.588 ;
        RECT 63.172 61.557 68.232 61.634 ;
        RECT 66.944 57.785 80 58.25 ;
        RECT 68.186 56.543 68.232 61.634 ;
        RECT 63.126 61.603 68.186 61.68 ;
        RECT 66.99 57.739 80 58.25 ;
        RECT 68.14 56.589 68.186 61.68 ;
        RECT 63.08 61.649 68.14 61.726 ;
        RECT 67.036 57.693 80 58.25 ;
        RECT 68.094 56.635 68.14 61.726 ;
        RECT 63.034 61.695 68.094 61.772 ;
        RECT 67.082 57.647 80 58.25 ;
        RECT 68.048 56.681 68.094 61.772 ;
        RECT 62.988 61.741 68.048 61.818 ;
        RECT 67.128 57.601 80 58.25 ;
        RECT 68.002 56.727 68.048 61.818 ;
        RECT 62.942 61.787 68.002 61.864 ;
        RECT 67.174 57.555 80 58.25 ;
        RECT 67.956 56.773 68.002 61.864 ;
        RECT 62.896 61.833 67.956 61.91 ;
        RECT 67.22 57.509 80 58.25 ;
        RECT 67.91 56.819 67.956 61.91 ;
        RECT 62.85 61.879 67.91 61.956 ;
        RECT 67.266 57.463 80 58.25 ;
        RECT 67.864 56.865 67.91 61.956 ;
        RECT 62.804 61.925 67.864 62.002 ;
        RECT 67.312 57.417 80 58.25 ;
        RECT 67.818 56.911 67.864 62.002 ;
        RECT 62.758 61.971 67.818 62.048 ;
        RECT 67.358 57.371 80 58.25 ;
        RECT 67.772 56.957 67.818 62.048 ;
        RECT 62.712 62.017 67.772 62.094 ;
        RECT 67.404 57.325 80 58.25 ;
        RECT 67.726 57.003 67.772 62.094 ;
        RECT 62.666 62.063 67.726 62.14 ;
        RECT 67.45 57.279 80 58.25 ;
        RECT 67.68 57.049 67.726 62.14 ;
        RECT 62.62 62.109 67.68 62.186 ;
        RECT 67.496 57.233 80 58.25 ;
        RECT 67.634 57.095 67.68 62.186 ;
        RECT 62.574 62.155 67.634 62.232 ;
        RECT 67.542 57.187 80 58.25 ;
        RECT 67.588 57.141 67.634 62.232 ;
        RECT 62.528 62.201 67.588 62.278 ;
        RECT 62.482 62.247 67.542 62.324 ;
        RECT 62.436 62.293 67.496 62.37 ;
        RECT 62.39 62.339 67.45 62.416 ;
        RECT 62.344 62.385 67.404 62.462 ;
        RECT 62.298 62.431 67.358 62.508 ;
        RECT 62.252 62.477 67.312 62.554 ;
        RECT 62.206 62.523 67.266 62.6 ;
        RECT 62.16 62.569 67.22 62.646 ;
        RECT 62.114 62.615 67.174 62.692 ;
        RECT 62.068 62.661 67.128 62.738 ;
        RECT 62.022 62.707 67.082 62.784 ;
        RECT 61.976 62.753 67.036 62.83 ;
        RECT 61.93 62.799 66.99 62.876 ;
        RECT 61.884 62.845 66.944 62.922 ;
        RECT 61.838 62.891 66.898 62.968 ;
        RECT 61.792 62.937 66.852 63.014 ;
        RECT 61.746 62.983 66.806 63.06 ;
        RECT 61.7 63.029 66.76 63.106 ;
        RECT 61.654 63.075 66.714 63.152 ;
        RECT 61.608 63.121 66.668 63.198 ;
        RECT 61.562 63.167 66.622 63.244 ;
        RECT 61.516 63.213 66.576 63.29 ;
        RECT 61.47 63.259 66.53 63.336 ;
        RECT 61.424 63.305 66.484 63.382 ;
        RECT 61.378 63.351 66.438 63.428 ;
        RECT 61.332 63.397 66.392 63.474 ;
        RECT 61.286 63.443 66.346 63.52 ;
        RECT 61.24 63.489 66.3 63.566 ;
        RECT 61.194 63.535 66.254 63.612 ;
        RECT 61.148 63.581 66.208 63.658 ;
        RECT 61.102 63.627 66.162 63.704 ;
        RECT 61.056 63.673 66.116 63.75 ;
        RECT 61.01 63.719 66.07 63.796 ;
        RECT 60.964 63.765 66.024 63.842 ;
        RECT 60.918 63.811 65.978 63.888 ;
        RECT 60.872 63.857 65.932 63.934 ;
        RECT 60.826 63.903 65.886 63.98 ;
        RECT 60.78 63.949 65.84 64.026 ;
        RECT 60.734 63.995 65.794 64.072 ;
        RECT 60.688 64.041 65.748 64.118 ;
        RECT 60.642 64.087 65.702 64.164 ;
        RECT 60.596 64.133 65.656 64.21 ;
        RECT 60.55 64.179 65.61 64.256 ;
        RECT 60.504 64.225 65.564 64.302 ;
        RECT 60.458 64.271 65.518 64.348 ;
        RECT 60.412 64.317 65.472 64.394 ;
        RECT 60.366 64.363 65.426 64.44 ;
        RECT 60.32 64.409 65.38 64.486 ;
        RECT 60.274 64.455 65.334 64.532 ;
        RECT 60.228 64.501 65.288 64.578 ;
        RECT 60.182 64.547 65.242 64.624 ;
        RECT 60.136 64.593 65.196 64.67 ;
        RECT 60.09 64.639 65.15 64.716 ;
        RECT 60.044 64.685 65.104 64.762 ;
        RECT 59.998 64.731 65.058 64.808 ;
        RECT 59.952 64.777 65.012 64.854 ;
        RECT 59.906 64.823 64.966 64.9 ;
        RECT 59.86 64.869 64.92 64.946 ;
        RECT 59.814 64.915 64.874 64.992 ;
        RECT 59.768 64.961 64.828 65.038 ;
        RECT 59.722 65.007 64.782 65.084 ;
        RECT 59.676 65.053 64.736 65.13 ;
        RECT 59.63 65.099 64.69 65.176 ;
        RECT 59.584 65.145 64.644 65.222 ;
        RECT 59.538 65.191 64.598 65.268 ;
        RECT 59.492 65.237 64.552 65.314 ;
        RECT 59.446 65.283 64.506 65.36 ;
        RECT 59.4 65.329 64.46 65.406 ;
        RECT 59.354 65.375 64.414 65.452 ;
        RECT 59.308 65.421 64.368 65.498 ;
        RECT 59.262 65.467 64.322 65.544 ;
        RECT 59.216 65.513 64.276 65.59 ;
        RECT 59.17 65.559 64.23 65.636 ;
        RECT 59.124 65.605 64.184 65.682 ;
        RECT 59.078 65.651 64.138 65.728 ;
        RECT 59.032 65.697 64.092 65.774 ;
        RECT 58.986 65.743 64.046 65.82 ;
        RECT 58.94 65.789 64 65.866 ;
        RECT 58.894 65.835 63.954 65.912 ;
        RECT 58.848 65.881 63.908 65.958 ;
        RECT 58.802 65.927 63.862 66.004 ;
        RECT 58.756 65.973 63.816 66.05 ;
        RECT 58.71 66.019 63.77 66.096 ;
        RECT 58.664 66.065 63.724 66.142 ;
        RECT 58.618 66.111 63.678 66.188 ;
        RECT 58.572 66.157 63.632 66.234 ;
        RECT 58.526 66.203 63.586 66.28 ;
        RECT 58.48 66.249 63.54 66.326 ;
        RECT 58.434 66.295 63.494 66.372 ;
        RECT 58.388 66.341 63.448 66.418 ;
        RECT 58.342 66.387 63.402 66.464 ;
        RECT 58.25 66.479 63.356 66.51 ;
        RECT 58.296 66.433 63.356 66.51 ;
        RECT 58.238 66.508 63.31 66.556 ;
        RECT 58.192 66.537 63.264 66.602 ;
        RECT 58.146 66.583 63.218 66.648 ;
        RECT 58.1 66.629 63.172 66.694 ;
        RECT 58.054 66.675 63.126 66.74 ;
        RECT 58.008 66.721 63.08 66.786 ;
        RECT 57.962 66.767 63.034 66.832 ;
        RECT 57.916 66.813 62.988 66.878 ;
        RECT 57.87 66.859 62.942 66.924 ;
        RECT 57.824 66.905 62.896 66.97 ;
        RECT 57.778 66.951 62.85 67.016 ;
        RECT 57.732 66.997 62.804 67.062 ;
        RECT 57.686 67.043 62.758 67.108 ;
        RECT 57.64 67.089 62.712 67.154 ;
        RECT 57.594 67.135 62.666 67.2 ;
        RECT 57.548 67.181 62.62 67.246 ;
        RECT 57.502 67.227 62.574 67.292 ;
        RECT 57.456 67.273 62.528 67.338 ;
        RECT 57.41 67.319 62.482 67.384 ;
        RECT 57.364 67.365 62.436 67.43 ;
        RECT 57.318 67.411 62.39 67.476 ;
        RECT 57.272 67.457 62.344 67.522 ;
        RECT 57.226 67.503 62.298 67.568 ;
        RECT 57.18 67.549 62.252 67.614 ;
        RECT 57.134 67.595 62.206 67.66 ;
        RECT 57.088 67.641 62.16 67.706 ;
        RECT 57.042 67.687 62.114 67.752 ;
        RECT 56.996 67.733 62.068 67.798 ;
        RECT 56.95 67.779 62.022 67.844 ;
        RECT 56.904 67.825 61.976 67.89 ;
        RECT 56.858 67.871 61.93 67.936 ;
        RECT 56.812 67.917 61.884 67.982 ;
        RECT 56.766 67.963 61.838 68.028 ;
        RECT 56.72 68.009 61.792 68.074 ;
        RECT 56.674 68.055 61.746 68.12 ;
        RECT 56.628 68.101 61.7 68.166 ;
        RECT 56.582 68.147 61.654 68.212 ;
        RECT 56.536 68.193 61.608 68.258 ;
        RECT 56.49 68.239 61.562 68.304 ;
        RECT 56.444 68.285 61.516 68.35 ;
        RECT 56.398 68.331 61.47 68.396 ;
        RECT 56.352 68.377 61.424 68.442 ;
        RECT 56.306 68.423 61.378 68.488 ;
        RECT 56.26 68.469 61.332 68.534 ;
        RECT 56.214 68.515 61.286 68.58 ;
        RECT 56.168 68.561 61.24 68.626 ;
        RECT 56.122 68.607 61.194 68.672 ;
        RECT 56.076 68.653 61.148 68.718 ;
        RECT 56.03 68.699 61.102 68.764 ;
        RECT 55.984 68.745 61.056 68.81 ;
        RECT 55.938 68.791 61.01 68.856 ;
        RECT 55.892 68.837 60.964 68.902 ;
        RECT 55.846 68.883 60.918 68.948 ;
        RECT 55.8 68.929 60.872 68.994 ;
        RECT 55.754 68.975 60.826 69.04 ;
        RECT 55.708 69.021 60.78 69.086 ;
        RECT 55.662 69.067 60.734 69.132 ;
        RECT 55.616 69.113 60.688 69.178 ;
        RECT 55.57 69.159 60.642 69.224 ;
        RECT 55.524 69.205 60.596 69.27 ;
        RECT 55.478 69.251 60.55 69.316 ;
        RECT 55.432 69.297 60.504 69.362 ;
        RECT 55.386 69.343 60.458 69.408 ;
        RECT 55.34 69.389 60.412 69.454 ;
        RECT 55.294 69.435 60.366 69.5 ;
        RECT 55.248 69.481 60.32 69.546 ;
        RECT 55.202 69.527 60.274 69.592 ;
        RECT 55.156 69.573 60.228 69.638 ;
        RECT 55.11 69.619 60.182 69.684 ;
        RECT 55.064 69.665 60.136 69.73 ;
        RECT 55.018 69.711 60.09 69.776 ;
        RECT 54.972 69.757 60.044 69.822 ;
        RECT 54.926 69.803 59.998 69.868 ;
        RECT 54.88 69.849 59.952 69.914 ;
        RECT 54.834 69.895 59.906 69.96 ;
        RECT 54.788 69.941 59.86 70.006 ;
        RECT 54.742 69.987 59.814 70.052 ;
        RECT 54.696 70.033 59.768 70.098 ;
        RECT 54.65 70.079 59.722 70.144 ;
        RECT 54.65 70.079 59.676 70.19 ;
        RECT 54.65 70.079 59.63 70.236 ;
        RECT 54.65 70.079 59.584 70.282 ;
        RECT 54.65 70.079 59.538 70.328 ;
        RECT 54.65 70.079 59.492 70.374 ;
        RECT 54.65 70.079 59.446 70.42 ;
        RECT 54.65 70.079 59.4 70.466 ;
        RECT 54.65 70.079 59.354 70.512 ;
        RECT 54.65 70.079 59.308 70.558 ;
        RECT 54.65 70.079 59.262 70.604 ;
        RECT 54.65 70.079 59.216 70.65 ;
        RECT 54.65 70.079 59.17 70.696 ;
        RECT 54.65 70.079 59.124 70.742 ;
        RECT 54.65 70.079 59.078 70.788 ;
        RECT 54.65 70.079 59.032 70.834 ;
        RECT 54.65 70.079 58.986 70.88 ;
        RECT 54.65 70.079 58.94 70.926 ;
        RECT 54.65 70.079 58.894 70.972 ;
        RECT 54.65 70.079 58.848 71.018 ;
        RECT 54.65 70.079 58.802 71.064 ;
        RECT 54.65 70.079 58.756 71.11 ;
        RECT 54.65 70.079 58.71 71.156 ;
        RECT 54.65 70.079 58.664 71.202 ;
        RECT 54.65 70.079 58.618 71.248 ;
        RECT 54.65 70.079 58.572 71.294 ;
        RECT 54.65 70.079 58.526 71.34 ;
        RECT 54.65 70.079 58.48 71.386 ;
        RECT 54.65 70.079 58.434 71.432 ;
        RECT 54.65 70.079 58.388 71.478 ;
        RECT 54.65 70.079 58.342 71.524 ;
        RECT 54.65 70.079 58.296 71.57 ;
        RECT 54.65 70.079 58.25 80 ;
        RECT 70.102 54.65 80 58.25 ;
        RECT 66.484 58.245 71.593 58.26 ;
        RECT 65.058 59.671 70.148 59.718 ;
        RECT 70.072 54.665 70.102 59.756 ;
        RECT 65.012 59.717 70.072 59.794 ;
        RECT 65.104 59.625 70.194 59.672 ;
        RECT 70.026 54.703 70.072 59.794 ;
        RECT 64.966 59.763 70.026 59.84 ;
        RECT 65.15 59.579 70.24 59.626 ;
        RECT 69.98 54.749 70.026 59.84 ;
        RECT 64.92 59.809 69.98 59.886 ;
        RECT 65.196 59.533 70.286 59.58 ;
        RECT 69.934 54.795 69.98 59.886 ;
        RECT 64.874 59.855 69.934 59.932 ;
        RECT 65.242 59.487 70.332 59.534 ;
        RECT 69.888 54.841 69.934 59.932 ;
        RECT 64.828 59.901 69.888 59.978 ;
        RECT 65.288 59.441 70.378 59.488 ;
        RECT 69.842 54.887 69.888 59.978 ;
        RECT 64.782 59.947 69.842 60.024 ;
        RECT 65.334 59.395 70.424 59.442 ;
        RECT 69.796 54.933 69.842 60.024 ;
        RECT 64.736 59.993 69.796 60.07 ;
        RECT 65.38 59.349 70.47 59.396 ;
        RECT 69.75 54.979 69.796 60.07 ;
        RECT 64.69 60.039 69.75 60.116 ;
        RECT 65.426 59.303 70.516 59.35 ;
        RECT 69.704 55.025 69.75 60.116 ;
        RECT 64.644 60.085 69.704 60.162 ;
        RECT 65.472 59.257 70.562 59.304 ;
        RECT 69.658 55.071 69.704 60.162 ;
        RECT 64.598 60.131 69.658 60.208 ;
        RECT 65.518 59.211 70.608 59.258 ;
        RECT 69.612 55.117 69.658 60.208 ;
        RECT 64.552 60.177 69.612 60.254 ;
        RECT 65.564 59.165 70.654 59.212 ;
        RECT 69.566 55.163 69.612 60.254 ;
        RECT 64.506 60.223 69.566 60.3 ;
        RECT 65.61 59.119 70.7 59.166 ;
        RECT 69.52 55.209 69.566 60.3 ;
        RECT 64.46 60.269 69.52 60.346 ;
        RECT 65.656 59.073 70.746 59.12 ;
        RECT 69.474 55.255 69.52 60.346 ;
        RECT 64.414 60.315 69.474 60.392 ;
        RECT 65.702 59.027 70.792 59.074 ;
        RECT 69.428 55.301 69.474 60.392 ;
        RECT 64.368 60.361 69.428 60.438 ;
        RECT 65.748 58.981 70.838 59.028 ;
        RECT 69.382 55.347 69.428 60.438 ;
        RECT 64.322 60.407 69.382 60.484 ;
        RECT 65.794 58.935 70.884 58.982 ;
        RECT 69.336 55.393 69.382 60.484 ;
        RECT 64.276 60.453 69.336 60.53 ;
        RECT 65.84 58.889 70.93 58.936 ;
        RECT 69.29 55.439 69.336 60.53 ;
        RECT 64.23 60.499 69.29 60.576 ;
        RECT 65.886 58.843 70.976 58.89 ;
        RECT 69.244 55.485 69.29 60.576 ;
        RECT 64.184 60.545 69.244 60.622 ;
        RECT 65.932 58.797 71.022 58.844 ;
        RECT 69.198 55.531 69.244 60.622 ;
        RECT 64.138 60.591 69.198 60.668 ;
        RECT 65.978 58.751 71.068 58.798 ;
        RECT 69.152 55.577 69.198 60.668 ;
        RECT 64.092 60.637 69.152 60.714 ;
        RECT 66.024 58.705 71.114 58.752 ;
        RECT 69.106 55.623 69.152 60.714 ;
        RECT 64.046 60.683 69.106 60.76 ;
        RECT 66.07 58.659 71.16 58.706 ;
        RECT 69.06 55.669 69.106 60.76 ;
        RECT 64 60.729 69.06 60.806 ;
        RECT 66.116 58.613 71.206 58.66 ;
        RECT 69.014 55.715 69.06 60.806 ;
        RECT 63.954 60.775 69.014 60.852 ;
        RECT 66.162 58.567 71.252 58.614 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 75.946 68.75 80 72.35 ;
        RECT 70.912 73.761 75.992 73.818 ;
        RECT 75.938 68.754 75.946 73.845 ;
        RECT 70.866 73.807 75.938 73.872 ;
        RECT 70.958 73.715 76.038 73.772 ;
        RECT 75.892 68.781 75.938 73.872 ;
        RECT 70.82 73.853 75.892 73.918 ;
        RECT 71.004 73.669 76.084 73.726 ;
        RECT 75.846 68.827 75.892 73.918 ;
        RECT 70.774 73.899 75.846 73.964 ;
        RECT 71.05 73.623 76.13 73.68 ;
        RECT 75.8 68.873 75.846 73.964 ;
        RECT 70.728 73.945 75.8 74.01 ;
        RECT 71.096 73.577 76.176 73.634 ;
        RECT 75.754 68.919 75.8 74.01 ;
        RECT 70.682 73.991 75.754 74.056 ;
        RECT 71.142 73.531 76.222 73.588 ;
        RECT 75.708 68.965 75.754 74.056 ;
        RECT 70.636 74.037 75.708 74.102 ;
        RECT 71.188 73.485 76.268 73.542 ;
        RECT 75.662 69.011 75.708 74.102 ;
        RECT 70.59 74.083 75.662 74.148 ;
        RECT 71.234 73.439 76.314 73.496 ;
        RECT 75.616 69.057 75.662 74.148 ;
        RECT 70.544 74.129 75.616 74.194 ;
        RECT 71.28 73.393 76.36 73.45 ;
        RECT 75.57 69.103 75.616 74.194 ;
        RECT 70.498 74.175 75.57 74.24 ;
        RECT 71.326 73.347 76.406 73.404 ;
        RECT 75.524 69.149 75.57 74.24 ;
        RECT 70.452 74.221 75.524 74.286 ;
        RECT 71.372 73.301 76.452 73.358 ;
        RECT 75.478 69.195 75.524 74.286 ;
        RECT 70.406 74.267 75.478 74.332 ;
        RECT 71.418 73.255 76.498 73.312 ;
        RECT 75.432 69.241 75.478 74.332 ;
        RECT 70.36 74.313 75.432 74.378 ;
        RECT 71.464 73.209 76.544 73.266 ;
        RECT 75.386 69.287 75.432 74.378 ;
        RECT 70.314 74.359 75.386 74.424 ;
        RECT 71.51 73.163 76.59 73.22 ;
        RECT 75.34 69.333 75.386 74.424 ;
        RECT 70.268 74.405 75.34 74.47 ;
        RECT 71.556 73.117 76.636 73.174 ;
        RECT 75.294 69.379 75.34 74.47 ;
        RECT 70.222 74.451 75.294 74.516 ;
        RECT 71.602 73.071 76.682 73.128 ;
        RECT 75.248 69.425 75.294 74.516 ;
        RECT 70.176 74.497 75.248 74.562 ;
        RECT 71.648 73.025 76.728 73.082 ;
        RECT 75.202 69.471 75.248 74.562 ;
        RECT 70.13 74.543 75.202 74.608 ;
        RECT 71.694 72.979 76.774 73.036 ;
        RECT 75.156 69.517 75.202 74.608 ;
        RECT 70.084 74.589 75.156 74.654 ;
        RECT 71.74 72.933 76.82 72.99 ;
        RECT 75.11 69.563 75.156 74.654 ;
        RECT 70.038 74.635 75.11 74.7 ;
        RECT 71.786 72.887 76.866 72.944 ;
        RECT 75.064 69.609 75.11 74.7 ;
        RECT 69.992 74.681 75.064 74.746 ;
        RECT 71.832 72.841 76.912 72.898 ;
        RECT 75.018 69.655 75.064 74.746 ;
        RECT 69.946 74.727 75.018 74.792 ;
        RECT 71.878 72.795 76.958 72.852 ;
        RECT 74.972 69.701 75.018 74.792 ;
        RECT 69.9 74.773 74.972 74.838 ;
        RECT 71.924 72.749 77.004 72.806 ;
        RECT 74.926 69.747 74.972 74.838 ;
        RECT 69.854 74.819 74.926 74.884 ;
        RECT 71.97 72.703 77.05 72.76 ;
        RECT 74.88 69.793 74.926 74.884 ;
        RECT 69.808 74.865 74.88 74.93 ;
        RECT 72.016 72.657 77.096 72.714 ;
        RECT 74.834 69.839 74.88 74.93 ;
        RECT 69.762 74.911 74.834 74.976 ;
        RECT 72.062 72.611 77.142 72.668 ;
        RECT 74.788 69.885 74.834 74.976 ;
        RECT 69.716 74.957 74.788 75.022 ;
        RECT 72.108 72.565 77.188 72.622 ;
        RECT 74.742 69.931 74.788 75.022 ;
        RECT 69.67 75.003 74.742 75.068 ;
        RECT 72.154 72.519 77.234 72.576 ;
        RECT 74.696 69.977 74.742 75.068 ;
        RECT 69.624 75.049 74.696 75.114 ;
        RECT 72.2 72.473 77.28 72.53 ;
        RECT 74.65 70.023 74.696 75.114 ;
        RECT 69.578 75.095 74.65 75.16 ;
        RECT 72.246 72.427 77.326 72.484 ;
        RECT 74.604 70.069 74.65 75.16 ;
        RECT 69.532 75.141 74.604 75.206 ;
        RECT 72.292 72.381 77.372 72.438 ;
        RECT 74.558 70.115 74.604 75.206 ;
        RECT 69.486 75.187 74.558 75.252 ;
        RECT 72.338 72.352 77.418 72.392 ;
        RECT 74.512 70.161 74.558 75.252 ;
        RECT 69.44 75.233 74.512 75.298 ;
        RECT 72.35 72.323 77.437 72.36 ;
        RECT 74.466 70.207 74.512 75.298 ;
        RECT 69.394 75.279 74.466 75.344 ;
        RECT 72.396 72.277 80 72.35 ;
        RECT 74.42 70.253 74.466 75.344 ;
        RECT 69.348 75.325 74.42 75.39 ;
        RECT 72.442 72.231 80 72.35 ;
        RECT 74.374 70.299 74.42 75.39 ;
        RECT 69.302 75.371 74.374 75.436 ;
        RECT 72.488 72.185 80 72.35 ;
        RECT 74.328 70.345 74.374 75.436 ;
        RECT 69.256 75.417 74.328 75.482 ;
        RECT 72.534 72.139 80 72.35 ;
        RECT 74.282 70.391 74.328 75.482 ;
        RECT 69.21 75.463 74.282 75.528 ;
        RECT 72.58 72.093 80 72.35 ;
        RECT 74.236 70.437 74.282 75.528 ;
        RECT 69.164 75.509 74.236 75.574 ;
        RECT 72.626 72.047 80 72.35 ;
        RECT 74.19 70.483 74.236 75.574 ;
        RECT 69.118 75.555 74.19 75.62 ;
        RECT 72.672 72.001 80 72.35 ;
        RECT 74.144 70.529 74.19 75.62 ;
        RECT 69.072 75.601 74.144 75.666 ;
        RECT 72.718 71.955 80 72.35 ;
        RECT 74.098 70.575 74.144 75.666 ;
        RECT 69.026 75.647 74.098 75.712 ;
        RECT 72.764 71.909 80 72.35 ;
        RECT 74.052 70.621 74.098 75.712 ;
        RECT 68.98 75.693 74.052 75.758 ;
        RECT 72.81 71.863 80 72.35 ;
        RECT 74.006 70.667 74.052 75.758 ;
        RECT 68.934 75.739 74.006 75.804 ;
        RECT 72.856 71.817 80 72.35 ;
        RECT 73.96 70.713 74.006 75.804 ;
        RECT 68.888 75.785 73.96 75.85 ;
        RECT 72.902 71.771 80 72.35 ;
        RECT 73.914 70.759 73.96 75.85 ;
        RECT 68.842 75.831 73.914 75.896 ;
        RECT 72.948 71.725 80 72.35 ;
        RECT 73.868 70.805 73.914 75.896 ;
        RECT 68.796 75.877 73.868 75.942 ;
        RECT 72.994 71.679 80 72.35 ;
        RECT 73.822 70.851 73.868 75.942 ;
        RECT 73.04 71.633 80 72.35 ;
        RECT 73.776 70.897 73.822 75.988 ;
        RECT 73.086 71.587 80 72.35 ;
        RECT 73.73 70.943 73.776 76.034 ;
        RECT 73.132 71.541 80 72.35 ;
        RECT 73.684 70.989 73.73 76.08 ;
        RECT 73.178 71.495 80 72.35 ;
        RECT 73.638 71.035 73.684 76.126 ;
        RECT 73.224 71.449 80 72.35 ;
        RECT 73.592 71.081 73.638 76.172 ;
        RECT 73.27 71.403 80 72.35 ;
        RECT 73.546 71.127 73.592 76.218 ;
        RECT 73.316 71.357 80 72.35 ;
        RECT 73.5 71.173 73.546 76.264 ;
        RECT 73.362 71.311 80 72.35 ;
        RECT 73.454 71.219 73.5 76.31 ;
        RECT 68.75 75.923 73.454 76.356 ;
        RECT 73.408 71.265 80 72.35 ;
        RECT 68.75 75.923 73.408 76.402 ;
        RECT 68.75 75.923 73.362 76.448 ;
        RECT 68.75 75.923 73.316 76.494 ;
        RECT 68.75 75.923 73.27 76.54 ;
        RECT 68.75 75.923 73.224 76.586 ;
        RECT 68.75 75.923 73.178 76.632 ;
        RECT 68.75 75.923 73.132 76.678 ;
        RECT 68.75 75.923 73.086 76.724 ;
        RECT 68.75 75.923 73.04 76.77 ;
        RECT 68.75 75.923 72.994 76.816 ;
        RECT 68.75 75.923 72.948 76.862 ;
        RECT 68.75 75.923 72.902 76.908 ;
        RECT 68.75 75.923 72.856 76.954 ;
        RECT 68.75 75.923 72.81 77 ;
        RECT 68.75 75.923 72.764 77.046 ;
        RECT 68.75 75.923 72.718 77.092 ;
        RECT 68.75 75.923 72.672 77.138 ;
        RECT 68.75 75.923 72.626 77.184 ;
        RECT 68.75 75.923 72.58 77.23 ;
        RECT 68.75 75.923 72.534 77.276 ;
        RECT 68.75 75.923 72.488 77.322 ;
        RECT 68.75 75.923 72.442 77.368 ;
        RECT 68.75 75.923 72.396 77.414 ;
        RECT 68.75 75.923 72.35 80 ;
    END
    PORT
      LAYER IB ;
        RECT 74.004 64.044 80 67.644 ;
        RECT 70.41 67.615 75.495 67.654 ;
        RECT 68.938 69.087 74.004 69.138 ;
        RECT 68.984 69.041 74.05 69.112 ;
        RECT 73.998 64.047 74.004 69.138 ;
        RECT 69.03 68.995 74.096 69.066 ;
        RECT 73.952 64.073 73.998 69.164 ;
        RECT 68.892 69.133 73.952 69.21 ;
        RECT 69.076 68.949 74.142 69.02 ;
        RECT 73.906 64.119 73.952 69.21 ;
        RECT 68.846 69.179 73.906 69.256 ;
        RECT 69.122 68.903 74.188 68.974 ;
        RECT 73.86 64.165 73.906 69.256 ;
        RECT 68.8 69.225 73.86 69.302 ;
        RECT 69.168 68.857 74.234 68.928 ;
        RECT 73.814 64.211 73.86 69.302 ;
        RECT 68.754 69.271 73.814 69.348 ;
        RECT 69.214 68.811 74.28 68.882 ;
        RECT 73.768 64.257 73.814 69.348 ;
        RECT 68.708 69.317 73.768 69.394 ;
        RECT 69.26 68.765 74.326 68.836 ;
        RECT 73.722 64.303 73.768 69.394 ;
        RECT 68.662 69.363 73.722 69.44 ;
        RECT 69.306 68.719 74.372 68.79 ;
        RECT 73.676 64.349 73.722 69.44 ;
        RECT 68.616 69.409 73.676 69.486 ;
        RECT 69.352 68.673 74.418 68.744 ;
        RECT 73.63 64.395 73.676 69.486 ;
        RECT 68.57 69.455 73.63 69.532 ;
        RECT 69.398 68.627 74.464 68.698 ;
        RECT 73.584 64.441 73.63 69.532 ;
        RECT 68.524 69.501 73.584 69.578 ;
        RECT 69.444 68.581 74.51 68.652 ;
        RECT 73.538 64.487 73.584 69.578 ;
        RECT 68.478 69.547 73.538 69.624 ;
        RECT 69.49 68.535 74.556 68.606 ;
        RECT 73.492 64.533 73.538 69.624 ;
        RECT 68.432 69.593 73.492 69.67 ;
        RECT 69.536 68.489 74.602 68.56 ;
        RECT 73.446 64.579 73.492 69.67 ;
        RECT 68.386 69.639 73.446 69.716 ;
        RECT 69.582 68.443 74.648 68.514 ;
        RECT 73.4 64.625 73.446 69.716 ;
        RECT 68.34 69.685 73.4 69.762 ;
        RECT 69.628 68.397 74.694 68.468 ;
        RECT 73.354 64.671 73.4 69.762 ;
        RECT 68.294 69.731 73.354 69.808 ;
        RECT 69.674 68.351 74.74 68.422 ;
        RECT 73.308 64.717 73.354 69.808 ;
        RECT 68.248 69.777 73.308 69.854 ;
        RECT 69.72 68.305 74.786 68.376 ;
        RECT 73.262 64.763 73.308 69.854 ;
        RECT 68.202 69.823 73.262 69.9 ;
        RECT 69.766 68.259 74.832 68.33 ;
        RECT 73.216 64.809 73.262 69.9 ;
        RECT 68.156 69.869 73.216 69.946 ;
        RECT 69.812 68.213 74.878 68.284 ;
        RECT 73.17 64.855 73.216 69.946 ;
        RECT 68.11 69.915 73.17 69.992 ;
        RECT 69.858 68.167 74.924 68.238 ;
        RECT 73.124 64.901 73.17 69.992 ;
        RECT 68.064 69.961 73.124 70.038 ;
        RECT 69.904 68.121 74.97 68.192 ;
        RECT 73.078 64.947 73.124 70.038 ;
        RECT 68.018 70.007 73.078 70.084 ;
        RECT 69.95 68.075 75.016 68.146 ;
        RECT 73.032 64.993 73.078 70.084 ;
        RECT 67.972 70.053 73.032 70.13 ;
        RECT 69.996 68.029 75.062 68.1 ;
        RECT 72.986 65.039 73.032 70.13 ;
        RECT 67.926 70.099 72.986 70.176 ;
        RECT 70.042 67.983 75.108 68.054 ;
        RECT 72.94 65.085 72.986 70.176 ;
        RECT 67.88 70.145 72.94 70.222 ;
        RECT 70.088 67.937 75.154 68.008 ;
        RECT 72.894 65.131 72.94 70.222 ;
        RECT 67.834 70.191 72.894 70.268 ;
        RECT 70.134 67.891 75.2 67.962 ;
        RECT 72.848 65.177 72.894 70.268 ;
        RECT 67.788 70.237 72.848 70.314 ;
        RECT 70.18 67.845 75.246 67.916 ;
        RECT 72.802 65.223 72.848 70.314 ;
        RECT 67.742 70.283 72.802 70.36 ;
        RECT 70.226 67.799 75.292 67.87 ;
        RECT 72.756 65.269 72.802 70.36 ;
        RECT 67.65 70.375 72.756 70.406 ;
        RECT 67.696 70.329 72.756 70.406 ;
        RECT 70.272 67.753 75.338 67.824 ;
        RECT 72.71 65.315 72.756 70.406 ;
        RECT 67.638 70.404 72.71 70.452 ;
        RECT 70.318 67.707 75.384 67.778 ;
        RECT 72.664 65.361 72.71 70.452 ;
        RECT 67.592 70.433 72.664 70.498 ;
        RECT 70.364 67.661 75.43 67.732 ;
        RECT 72.618 65.407 72.664 70.498 ;
        RECT 67.546 70.479 72.618 70.544 ;
        RECT 70.41 67.615 75.476 67.686 ;
        RECT 72.572 65.453 72.618 70.544 ;
        RECT 67.5 70.525 72.572 70.59 ;
        RECT 70.456 67.569 80 67.644 ;
        RECT 72.526 65.499 72.572 70.59 ;
        RECT 67.454 70.571 72.526 70.636 ;
        RECT 70.502 67.523 80 67.644 ;
        RECT 72.48 65.545 72.526 70.636 ;
        RECT 67.408 70.617 72.48 70.682 ;
        RECT 70.548 67.477 80 67.644 ;
        RECT 72.434 65.591 72.48 70.682 ;
        RECT 67.362 70.663 72.434 70.728 ;
        RECT 70.594 67.431 80 67.644 ;
        RECT 72.388 65.637 72.434 70.728 ;
        RECT 67.316 70.709 72.388 70.774 ;
        RECT 70.64 67.385 80 67.644 ;
        RECT 72.342 65.683 72.388 70.774 ;
        RECT 67.27 70.755 72.342 70.82 ;
        RECT 70.686 67.339 80 67.644 ;
        RECT 72.296 65.729 72.342 70.82 ;
        RECT 67.224 70.801 72.296 70.866 ;
        RECT 70.732 67.293 80 67.644 ;
        RECT 72.25 65.775 72.296 70.866 ;
        RECT 67.178 70.847 72.25 70.912 ;
        RECT 70.778 67.247 80 67.644 ;
        RECT 72.204 65.821 72.25 70.912 ;
        RECT 67.132 70.893 72.204 70.958 ;
        RECT 70.824 67.201 80 67.644 ;
        RECT 72.158 65.867 72.204 70.958 ;
        RECT 67.086 70.939 72.158 71.004 ;
        RECT 70.87 67.155 80 67.644 ;
        RECT 72.112 65.913 72.158 71.004 ;
        RECT 67.04 70.985 72.112 71.05 ;
        RECT 70.916 67.109 80 67.644 ;
        RECT 72.066 65.959 72.112 71.05 ;
        RECT 66.994 71.031 72.066 71.096 ;
        RECT 70.962 67.063 80 67.644 ;
        RECT 72.02 66.005 72.066 71.096 ;
        RECT 66.948 71.077 72.02 71.142 ;
        RECT 71.008 67.017 80 67.644 ;
        RECT 71.974 66.051 72.02 71.142 ;
        RECT 66.902 71.123 71.974 71.188 ;
        RECT 71.054 66.971 80 67.644 ;
        RECT 71.928 66.097 71.974 71.188 ;
        RECT 66.856 71.169 71.928 71.234 ;
        RECT 71.1 66.925 80 67.644 ;
        RECT 71.882 66.143 71.928 71.234 ;
        RECT 66.81 71.215 71.882 71.28 ;
        RECT 71.146 66.879 80 67.644 ;
        RECT 71.836 66.189 71.882 71.28 ;
        RECT 66.764 71.261 71.836 71.326 ;
        RECT 71.192 66.833 80 67.644 ;
        RECT 71.79 66.235 71.836 71.326 ;
        RECT 66.718 71.307 71.79 71.372 ;
        RECT 71.238 66.787 80 67.644 ;
        RECT 71.744 66.281 71.79 71.372 ;
        RECT 66.672 71.353 71.744 71.418 ;
        RECT 71.284 66.741 80 67.644 ;
        RECT 71.698 66.327 71.744 71.418 ;
        RECT 66.626 71.399 71.698 71.464 ;
        RECT 71.33 66.695 80 67.644 ;
        RECT 71.652 66.373 71.698 71.464 ;
        RECT 66.58 71.445 71.652 71.51 ;
        RECT 71.376 66.649 80 67.644 ;
        RECT 71.606 66.419 71.652 71.51 ;
        RECT 66.534 71.491 71.606 71.556 ;
        RECT 71.422 66.603 80 67.644 ;
        RECT 71.56 66.465 71.606 71.556 ;
        RECT 66.488 71.537 71.56 71.602 ;
        RECT 71.468 66.557 80 67.644 ;
        RECT 71.514 66.511 71.56 71.602 ;
        RECT 66.442 71.583 71.514 71.648 ;
        RECT 66.396 71.629 71.468 71.694 ;
        RECT 66.35 71.675 71.422 71.74 ;
        RECT 66.304 71.721 71.376 71.786 ;
        RECT 66.258 71.767 71.33 71.832 ;
        RECT 66.212 71.813 71.284 71.878 ;
        RECT 66.166 71.859 71.238 71.924 ;
        RECT 66.12 71.905 71.192 71.97 ;
        RECT 66.074 71.951 71.146 72.016 ;
        RECT 66.028 71.997 71.1 72.062 ;
        RECT 65.982 72.043 71.054 72.108 ;
        RECT 65.936 72.089 71.008 72.154 ;
        RECT 65.89 72.135 70.962 72.2 ;
        RECT 65.844 72.181 70.916 72.246 ;
        RECT 65.798 72.227 70.87 72.292 ;
        RECT 65.752 72.273 70.824 72.338 ;
        RECT 65.706 72.319 70.778 72.384 ;
        RECT 65.66 72.365 70.732 72.43 ;
        RECT 65.614 72.411 70.686 72.476 ;
        RECT 65.568 72.457 70.64 72.522 ;
        RECT 65.522 72.503 70.594 72.568 ;
        RECT 65.476 72.549 70.548 72.614 ;
        RECT 65.43 72.595 70.502 72.66 ;
        RECT 65.384 72.641 70.456 72.706 ;
        RECT 65.338 72.687 70.41 72.752 ;
        RECT 65.292 72.733 70.364 72.798 ;
        RECT 65.246 72.779 70.318 72.844 ;
        RECT 65.2 72.825 70.272 72.89 ;
        RECT 65.154 72.871 70.226 72.936 ;
        RECT 65.108 72.917 70.18 72.982 ;
        RECT 65.062 72.963 70.134 73.028 ;
        RECT 65.016 73.009 70.088 73.074 ;
        RECT 64.97 73.055 70.042 73.12 ;
        RECT 64.924 73.101 69.996 73.166 ;
        RECT 64.878 73.147 69.95 73.212 ;
        RECT 64.832 73.193 69.904 73.258 ;
        RECT 64.786 73.239 69.858 73.304 ;
        RECT 64.74 73.285 69.812 73.35 ;
        RECT 64.694 73.331 69.766 73.396 ;
        RECT 64.648 73.377 69.72 73.442 ;
        RECT 64.602 73.423 69.674 73.488 ;
        RECT 64.556 73.469 69.628 73.534 ;
        RECT 64.51 73.515 69.582 73.58 ;
        RECT 64.464 73.561 69.536 73.626 ;
        RECT 64.418 73.607 69.49 73.672 ;
        RECT 64.372 73.653 69.444 73.718 ;
        RECT 64.326 73.699 69.398 73.764 ;
        RECT 64.28 73.745 69.352 73.81 ;
        RECT 64.234 73.791 69.306 73.856 ;
        RECT 64.188 73.837 69.26 73.902 ;
        RECT 64.142 73.883 69.214 73.948 ;
        RECT 64.096 73.929 69.168 73.994 ;
        RECT 64.05 73.975 69.122 74.04 ;
        RECT 64.05 73.975 69.076 74.086 ;
        RECT 64.05 73.975 69.03 74.132 ;
        RECT 64.05 73.975 68.984 74.178 ;
        RECT 64.05 73.975 68.938 74.224 ;
        RECT 64.05 73.975 68.892 74.27 ;
        RECT 64.05 73.975 68.846 74.316 ;
        RECT 64.05 73.975 68.8 74.362 ;
        RECT 64.05 73.975 68.754 74.408 ;
        RECT 64.05 73.975 68.708 74.454 ;
        RECT 64.05 73.975 68.662 74.5 ;
        RECT 64.05 73.975 68.616 74.546 ;
        RECT 64.05 73.975 68.57 74.592 ;
        RECT 64.05 73.975 68.524 74.638 ;
        RECT 64.05 73.975 68.478 74.684 ;
        RECT 64.05 73.975 68.432 74.73 ;
        RECT 64.05 73.975 68.386 74.776 ;
        RECT 64.05 73.975 68.34 74.822 ;
        RECT 64.05 73.975 68.294 74.868 ;
        RECT 64.05 73.975 68.248 74.914 ;
        RECT 64.05 73.975 68.202 74.96 ;
        RECT 64.05 73.975 68.156 75.006 ;
        RECT 64.05 73.975 68.11 75.052 ;
        RECT 64.05 73.975 68.064 75.098 ;
        RECT 64.05 73.975 68.018 75.144 ;
        RECT 64.05 73.975 67.972 75.19 ;
        RECT 64.05 73.975 67.926 75.236 ;
        RECT 64.05 73.975 67.88 75.282 ;
        RECT 64.05 73.975 67.834 75.328 ;
        RECT 64.05 73.975 67.788 75.374 ;
        RECT 64.05 73.975 67.742 75.42 ;
        RECT 64.05 73.975 67.696 75.466 ;
        RECT 64.05 73.975 67.65 80 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 80 ;
    LAYER M1 ;
      RECT 0 0 80 80 ;
    LAYER V1 ;
      RECT 0 0 80 80 ;
    LAYER M2 ;
      RECT 0 0 80 80 ;
    LAYER A1 ;
      RECT 0 0 80 80 ;
    LAYER C2 ;
      RECT 0 0 80 80 ;
    LAYER IA ;
      RECT 0 0 80 80 ;
    LAYER XA ;
      RECT 0 0 80 80 ;
    LAYER YX ;
      RECT 0 0 80 80 ;
    LAYER IB ;
      RECT 0 0 80 80 ;
    LAYER CB ;
      RECT 0 0 80 80 ;
    LAYER AY ;
      RECT 0 0 80 80 ;
    LAYER C1 ;
      RECT 0 0 80 80 ;
    LAYER C5 ;
      RECT 0 0 80 80 ;
    LAYER C4 ;
      RECT 0 0 80 80 ;
    LAYER C3 ;
      RECT 0 0 80 80 ;
    LAYER A5 ;
      RECT 0 0 80 80 ;
    LAYER A4 ;
      RECT 0 0 80 80 ;
    LAYER A3 ;
      RECT 0 0 80 80 ;
    LAYER A2 ;
      RECT 0 0 80 80 ;
    LAYER C6 ;
      RECT 0 0 80 80 ;
  END
END RIIO_EG1D80V_CORNER_45

MACRO RIIO_EG1D80V_CORNER_EG
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CORNER_EG 0 0 ;
  SIZE 80 BY 80 ;
  SYMMETRY X Y ;
  SITE corner_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 1.85 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 68.75 1.85 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 1.85 67.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 1.85 62.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 54.65 1.85 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.95 1.85 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 1.85 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 1.85 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 1.85 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 1.85 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 1.85 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 21.75 1.85 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 1.85 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 1.85 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 1.85 11.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 2.95 1.85 6.55 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 54.65 80 58.25 ;
        RECT 54.65 54.65 58.25 80 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 45.25 80 48.85 ;
        RECT 45.25 45.25 48.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 40.55 80 44.15 ;
        RECT 40.55 40.55 44.15 80 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 26.45 80 30.05 ;
        RECT 26.45 26.45 30.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 17.05 80 20.65 ;
        RECT 17.05 17.05 20.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 3.67 3.67 80 6.55 ;
        RECT 3.67 3.67 6.55 80 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 2.95 0 6.55 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 0 25.35 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 49.95 80 53.55 ;
        RECT 49.95 49.95 53.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 35.85 80 39.45 ;
        RECT 35.85 35.85 39.45 80 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 31.15 80 34.75 ;
        RECT 31.15 31.15 34.75 80 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 12.35 80 15.95 ;
        RECT 12.35 12.35 15.95 80 ;
    END
    PORT
      LAYER IB ;
        RECT 7.65 7.65 80 11.25 ;
        RECT 7.65 7.65 11.25 80 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 68.75 68.75 80 72.35 ;
        RECT 68.75 68.75 72.35 80 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 64.05 80 67.65 ;
        RECT 64.05 64.05 67.65 80 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 73.45 73.45 80 77.05 ;
        RECT 73.45 73.45 77.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 59.35 80 62.95 ;
        RECT 59.35 59.35 62.95 80 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 80 ;
    LAYER M1 ;
      RECT 0 0 80 80 ;
    LAYER V1 ;
      RECT 0 0 80 80 ;
    LAYER M2 ;
      RECT 0 0 80 80 ;
    LAYER A1 ;
      RECT 0 0 80 80 ;
    LAYER C2 ;
      RECT 0 0 80 80 ;
    LAYER IA ;
      RECT 0 0 80 80 ;
    LAYER XA ;
      RECT 0 0 80 80 ;
    LAYER YX ;
      RECT 0 0 80 80 ;
    LAYER IB ;
      RECT 0 0 80 80 ;
    LAYER CB ;
      RECT 0 0 80 80 ;
    LAYER AY ;
      RECT 0 0 80 80 ;
    LAYER C1 ;
      RECT 0 0 80 80 ;
    LAYER C5 ;
      RECT 0 0 80 80 ;
    LAYER C4 ;
      RECT 0 0 80 80 ;
    LAYER C3 ;
      RECT 0 0 80 80 ;
    LAYER A5 ;
      RECT 0 0 80 80 ;
    LAYER A4 ;
      RECT 0 0 80 80 ;
    LAYER A3 ;
      RECT 0 0 80 80 ;
    LAYER A2 ;
      RECT 0 0 80 80 ;
    LAYER C6 ;
      RECT 0 0 80 80 ;
  END
END RIIO_EG1D80V_CORNER_EG

MACRO RIIO_EG1D80V_CORNER_HVT
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CORNER_HVT 0 0 ;
  SIZE 80 BY 80 ;
  SYMMETRY X Y ;
  SITE corner_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 1.85 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 68.75 1.85 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 1.85 67.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 1.85 62.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 54.65 1.85 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.95 1.85 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 1.85 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 1.85 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 1.85 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 1.85 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 1.85 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 21.75 1.85 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 1.85 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 1.85 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 1.85 11.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 2.95 1.85 6.55 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 54.65 80 58.25 ;
        RECT 54.65 54.65 58.25 80 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 45.25 80 48.85 ;
        RECT 45.25 45.25 48.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 40.55 80 44.15 ;
        RECT 40.55 40.55 44.15 80 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 26.45 80 30.05 ;
        RECT 26.45 26.45 30.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 17.05 80 20.65 ;
        RECT 17.05 17.05 20.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 3.67 3.67 80 6.55 ;
        RECT 3.67 3.67 6.55 80 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 2.95 0 6.55 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 0 25.35 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 49.95 80 53.55 ;
        RECT 49.95 49.95 53.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 35.85 80 39.45 ;
        RECT 35.85 35.85 39.45 80 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 31.15 80 34.75 ;
        RECT 31.15 31.15 34.75 80 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 12.35 80 15.95 ;
        RECT 12.35 12.35 15.95 80 ;
    END
    PORT
      LAYER IB ;
        RECT 7.65 7.65 80 11.25 ;
        RECT 7.65 7.65 11.25 80 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 68.75 68.75 80 72.35 ;
        RECT 68.75 68.75 72.35 80 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 64.05 80 67.65 ;
        RECT 64.05 64.05 67.65 80 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 73.45 73.45 80 77.05 ;
        RECT 73.45 73.45 77.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 59.35 80 62.95 ;
        RECT 59.35 59.35 62.95 80 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 80 ;
    LAYER M1 ;
      RECT 0 0 80 80 ;
    LAYER V1 ;
      RECT 0 0 80 80 ;
    LAYER M2 ;
      RECT 0 0 80 80 ;
    LAYER A1 ;
      RECT 0 0 80 80 ;
    LAYER C2 ;
      RECT 0 0 80 80 ;
    LAYER IA ;
      RECT 0 0 80 80 ;
    LAYER XA ;
      RECT 0 0 80 80 ;
    LAYER YX ;
      RECT 0 0 80 80 ;
    LAYER IB ;
      RECT 0 0 80 80 ;
    LAYER CB ;
      RECT 0 0 80 80 ;
    LAYER AY ;
      RECT 0 0 80 80 ;
    LAYER C1 ;
      RECT 0 0 80 80 ;
    LAYER C5 ;
      RECT 0 0 80 80 ;
    LAYER C4 ;
      RECT 0 0 80 80 ;
    LAYER C3 ;
      RECT 0 0 80 80 ;
    LAYER A5 ;
      RECT 0 0 80 80 ;
    LAYER A4 ;
      RECT 0 0 80 80 ;
    LAYER A3 ;
      RECT 0 0 80 80 ;
    LAYER A2 ;
      RECT 0 0 80 80 ;
    LAYER C6 ;
      RECT 0 0 80 80 ;
  END
END RIIO_EG1D80V_CORNER_HVT

MACRO RIIO_EG1D80V_CORNER_RVT
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CORNER_RVT 0 0 ;
  SIZE 80 BY 80 ;
  SYMMETRY X Y ;
  SITE corner_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 1.85 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 68.75 1.85 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 1.85 67.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 1.85 62.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 54.65 1.85 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.95 1.85 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 1.85 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 1.85 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 1.85 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 1.85 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 1.85 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 21.75 1.85 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 1.85 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 1.85 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 1.85 11.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 2.95 1.85 6.55 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 54.65 80 58.25 ;
        RECT 54.65 54.65 58.25 80 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 45.25 80 48.85 ;
        RECT 45.25 45.25 48.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 40.55 80 44.15 ;
        RECT 40.55 40.55 44.15 80 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 26.45 80 30.05 ;
        RECT 26.45 26.45 30.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 17.05 80 20.65 ;
        RECT 17.05 17.05 20.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 3.67 3.67 80 6.55 ;
        RECT 3.67 3.67 6.55 80 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 2.95 0 6.55 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 0 25.35 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 49.95 80 53.55 ;
        RECT 49.95 49.95 53.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 35.85 80 39.45 ;
        RECT 35.85 35.85 39.45 80 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 31.15 80 34.75 ;
        RECT 31.15 31.15 34.75 80 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 12.35 80 15.95 ;
        RECT 12.35 12.35 15.95 80 ;
    END
    PORT
      LAYER IB ;
        RECT 7.65 7.65 80 11.25 ;
        RECT 7.65 7.65 11.25 80 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 68.75 68.75 80 72.35 ;
        RECT 68.75 68.75 72.35 80 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 64.05 80 67.65 ;
        RECT 64.05 64.05 67.65 80 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 73.45 73.45 80 77.05 ;
        RECT 73.45 73.45 77.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 59.35 80 62.95 ;
        RECT 59.35 59.35 62.95 80 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 80 ;
    LAYER M1 ;
      RECT 0 0 80 80 ;
    LAYER V1 ;
      RECT 0 0 80 80 ;
    LAYER M2 ;
      RECT 0 0 80 80 ;
    LAYER A1 ;
      RECT 0 0 80 80 ;
    LAYER C2 ;
      RECT 0 0 80 80 ;
    LAYER IA ;
      RECT 0 0 80 80 ;
    LAYER XA ;
      RECT 0 0 80 80 ;
    LAYER YX ;
      RECT 0 0 80 80 ;
    LAYER IB ;
      RECT 0 0 80 80 ;
    LAYER CB ;
      RECT 0 0 80 80 ;
    LAYER AY ;
      RECT 0 0 80 80 ;
    LAYER C1 ;
      RECT 0 0 80 80 ;
    LAYER C5 ;
      RECT 0 0 80 80 ;
    LAYER C4 ;
      RECT 0 0 80 80 ;
    LAYER C3 ;
      RECT 0 0 80 80 ;
    LAYER A5 ;
      RECT 0 0 80 80 ;
    LAYER A4 ;
      RECT 0 0 80 80 ;
    LAYER A3 ;
      RECT 0 0 80 80 ;
    LAYER A2 ;
      RECT 0 0 80 80 ;
    LAYER C6 ;
      RECT 0 0 80 80 ;
  END
END RIIO_EG1D80V_CORNER_RVT

MACRO RIIO_EG1D80V_ANACORE_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ANACORE_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VESD3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 63.22955 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 7.36 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 52.45 78.15 52.95 80 ;
        RECT 51.675 78.15 52.175 80 ;
        RECT 50.9 78.15 51.4 80 ;
        RECT 50.125 78.15 50.625 80 ;
        RECT 49.35 78.15 49.85 80 ;
      LAYER M2 ;
        RECT 52.45 78.15 52.95 80 ;
        RECT 51.675 78.15 52.175 80 ;
        RECT 50.9 78.15 51.4 80 ;
        RECT 50.125 78.15 50.625 80 ;
        RECT 49.35 78.15 49.85 80 ;
      LAYER C1 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IA ;
        RECT 49.65 77.975 52.65 80 ;
    END
  END VESD3_B
  PIN VRES1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 75.6725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 19.55 78.15 20.05 80 ;
        RECT 18.775 78.15 19.275 80 ;
        RECT 18 78.15 18.5 80 ;
        RECT 17.225 78.15 17.725 80 ;
        RECT 16.45 78.15 16.95 80 ;
      LAYER M2 ;
        RECT 19.55 78.15 20.05 80 ;
        RECT 18.775 78.15 19.275 80 ;
        RECT 18 78.15 18.5 80 ;
        RECT 17.225 78.15 17.725 80 ;
        RECT 16.45 78.15 16.95 80 ;
      LAYER C1 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IA ;
        RECT 16.75 77.975 19.75 80 ;
    END
  END VRES1_B
  PIN VRES0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 72.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 16.735 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.4675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 14.85 78.15 15.35 80 ;
        RECT 14.075 78.15 14.575 80 ;
        RECT 13.3 78.15 13.8 80 ;
        RECT 12.525 78.15 13.025 80 ;
        RECT 11.75 78.15 12.25 80 ;
      LAYER M2 ;
        RECT 14.85 78.15 15.35 80 ;
        RECT 14.075 78.15 14.575 80 ;
        RECT 13.3 78.15 13.8 80 ;
        RECT 12.525 78.15 13.025 80 ;
        RECT 11.75 78.15 12.25 80 ;
      LAYER C1 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IA ;
        RECT 12.05 77.975 15.05 80 ;
    END
  END VRES0_B
  PIN VRES3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 72.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.4675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 47.75 78.15 48.25 80 ;
        RECT 46.975 78.15 47.475 80 ;
        RECT 46.2 78.15 46.7 80 ;
        RECT 45.425 78.15 45.925 80 ;
        RECT 44.65 78.15 45.15 80 ;
      LAYER M2 ;
        RECT 47.75 78.15 48.25 80 ;
        RECT 46.975 78.15 47.475 80 ;
        RECT 46.2 78.15 46.7 80 ;
        RECT 45.425 78.15 45.925 80 ;
        RECT 44.65 78.15 45.15 80 ;
      LAYER C1 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IA ;
        RECT 44.95 77.975 47.95 80 ;
    END
  END VRES3_B
  PIN VESD1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 24.25 78.15 24.75 80 ;
        RECT 23.475 78.15 23.975 80 ;
        RECT 22.7 78.15 23.2 80 ;
        RECT 21.925 78.15 22.425 80 ;
        RECT 21.15 78.15 21.65 80 ;
      LAYER M2 ;
        RECT 24.25 78.15 24.75 80 ;
        RECT 23.475 78.15 23.975 80 ;
        RECT 22.7 78.15 23.2 80 ;
        RECT 21.925 78.15 22.425 80 ;
        RECT 21.15 78.15 21.65 80 ;
      LAYER C1 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IA ;
        RECT 21.45 77.975 24.45 80 ;
    END
  END VESD1_B
  PIN VRES2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 75.6725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 7.36 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 43.05 78.15 43.55 80 ;
        RECT 42.275 78.15 42.775 80 ;
        RECT 41.5 78.15 42 80 ;
        RECT 40.725 78.15 41.225 80 ;
        RECT 39.95 78.15 40.45 80 ;
      LAYER M2 ;
        RECT 43.05 78.15 43.55 80 ;
        RECT 42.275 78.15 42.775 80 ;
        RECT 41.5 78.15 42 80 ;
        RECT 40.725 78.15 41.225 80 ;
        RECT 39.95 78.15 40.45 80 ;
      LAYER C1 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IA ;
        RECT 40.25 77.975 43.25 80 ;
    END
  END VRES2_B
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VESD0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 7.36 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 10.15 78.15 10.65 80 ;
        RECT 9.375 78.15 9.875 80 ;
        RECT 8.6 78.15 9.1 80 ;
        RECT 7.825 78.15 8.325 80 ;
        RECT 7.05 78.15 7.55 80 ;
      LAYER M2 ;
        RECT 10.15 78.15 10.65 80 ;
        RECT 9.375 78.15 9.875 80 ;
        RECT 8.6 78.15 9.1 80 ;
        RECT 7.825 78.15 8.325 80 ;
        RECT 7.05 78.15 7.55 80 ;
      LAYER C1 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IA ;
        RECT 7.35 77.975 10.35 80 ;
    END
  END VESD0_B
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 116.6975 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 493.9475 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 95.645 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 337.235 LAYER IA ;
    ANTENNAPARTIALMETALAREA 294.725 LAYER IB ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 12.59712 LAYER YX ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER XA ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A2 ;
    ANTENNADIFFAREA 150.1 LAYER C5 ;
    ANTENNADIFFAREA 150.1 LAYER C4 ;
    ANTENNADIFFAREA 150.1 LAYER C6 ;
    ANTENNADIFFAREA 150.1 LAYER IA ;
    ANTENNADIFFAREA 150.1 LAYER IB ;
    ANTENNADIFFAREA 150.1 LAYER C3 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 2.35 21.75 57.65 25.35 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN VESD2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 38.35 78.15 38.85 80 ;
        RECT 37.575 78.15 38.075 80 ;
        RECT 36.8 78.15 37.3 80 ;
        RECT 36.025 78.15 36.525 80 ;
        RECT 35.25 78.15 35.75 80 ;
      LAYER M2 ;
        RECT 38.35 78.15 38.85 80 ;
        RECT 37.575 78.15 38.075 80 ;
        RECT 36.8 78.15 37.3 80 ;
        RECT 36.025 78.15 36.525 80 ;
        RECT 35.25 78.15 35.75 80 ;
      LAYER C1 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IA ;
        RECT 35.55 77.975 38.55 80 ;
    END
  END VESD2_B
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_ANACORE_V

MACRO RIIO_EG1D80V_ANAIO_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ANAIO_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VESD3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 63.22955 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 7.36 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 52.45 78.15 52.95 80 ;
        RECT 51.675 78.15 52.175 80 ;
        RECT 50.9 78.15 51.4 80 ;
        RECT 50.125 78.15 50.625 80 ;
        RECT 49.35 78.15 49.85 80 ;
      LAYER M2 ;
        RECT 52.45 78.15 52.95 80 ;
        RECT 51.675 78.15 52.175 80 ;
        RECT 50.9 78.15 51.4 80 ;
        RECT 50.125 78.15 50.625 80 ;
        RECT 49.35 78.15 49.85 80 ;
      LAYER C1 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IA ;
        RECT 49.65 77.975 52.65 80 ;
    END
  END VESD3_B
  PIN VRES1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 75.6725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 19.55 78.15 20.05 80 ;
        RECT 18.775 78.15 19.275 80 ;
        RECT 18 78.15 18.5 80 ;
        RECT 17.225 78.15 17.725 80 ;
        RECT 16.45 78.15 16.95 80 ;
      LAYER M2 ;
        RECT 19.55 78.15 20.05 80 ;
        RECT 18.775 78.15 19.275 80 ;
        RECT 18 78.15 18.5 80 ;
        RECT 17.225 78.15 17.725 80 ;
        RECT 16.45 78.15 16.95 80 ;
      LAYER C1 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IA ;
        RECT 16.75 77.975 19.75 80 ;
    END
  END VRES1_B
  PIN VRES0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 72.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 16.735 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.4675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 14.85 78.15 15.35 80 ;
        RECT 14.075 78.15 14.575 80 ;
        RECT 13.3 78.15 13.8 80 ;
        RECT 12.525 78.15 13.025 80 ;
        RECT 11.75 78.15 12.25 80 ;
      LAYER M2 ;
        RECT 14.85 78.15 15.35 80 ;
        RECT 14.075 78.15 14.575 80 ;
        RECT 13.3 78.15 13.8 80 ;
        RECT 12.525 78.15 13.025 80 ;
        RECT 11.75 78.15 12.25 80 ;
      LAYER C1 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IA ;
        RECT 12.05 77.975 15.05 80 ;
    END
  END VRES0_B
  PIN VRES3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 72.8425 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 16.735 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.4675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 47.75 78.15 48.25 80 ;
        RECT 46.975 78.15 47.475 80 ;
        RECT 46.2 78.15 46.7 80 ;
        RECT 45.425 78.15 45.925 80 ;
        RECT 44.65 78.15 45.15 80 ;
      LAYER M2 ;
        RECT 47.75 78.15 48.25 80 ;
        RECT 46.975 78.15 47.475 80 ;
        RECT 46.2 78.15 46.7 80 ;
        RECT 45.425 78.15 45.925 80 ;
        RECT 44.65 78.15 45.15 80 ;
      LAYER C1 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IA ;
        RECT 44.95 77.975 47.95 80 ;
    END
  END VRES3_B
  PIN VESD1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 24.25 78.15 24.75 80 ;
        RECT 23.475 78.15 23.975 80 ;
        RECT 22.7 78.15 23.2 80 ;
        RECT 21.925 78.15 22.425 80 ;
        RECT 21.15 78.15 21.65 80 ;
      LAYER M2 ;
        RECT 24.25 78.15 24.75 80 ;
        RECT 23.475 78.15 23.975 80 ;
        RECT 22.7 78.15 23.2 80 ;
        RECT 21.925 78.15 22.425 80 ;
        RECT 21.15 78.15 21.65 80 ;
      LAYER C1 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IA ;
        RECT 21.45 77.975 24.45 80 ;
    END
  END VESD1_B
  PIN VRES2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 75.6725 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 7.36 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 43.05 78.15 43.55 80 ;
        RECT 42.275 78.15 42.775 80 ;
        RECT 41.5 78.15 42 80 ;
        RECT 40.725 78.15 41.225 80 ;
        RECT 39.95 78.15 40.45 80 ;
      LAYER M2 ;
        RECT 43.05 78.15 43.55 80 ;
        RECT 42.275 78.15 42.775 80 ;
        RECT 41.5 78.15 42 80 ;
        RECT 40.725 78.15 41.225 80 ;
        RECT 39.95 78.15 40.45 80 ;
      LAYER C1 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IA ;
        RECT 40.25 77.975 43.25 80 ;
    END
  END VRES2_B
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VESD0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 7.36 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 10.15 78.15 10.65 80 ;
        RECT 9.375 78.15 9.875 80 ;
        RECT 8.6 78.15 9.1 80 ;
        RECT 7.825 78.15 8.325 80 ;
        RECT 7.05 78.15 7.55 80 ;
      LAYER M2 ;
        RECT 10.15 78.15 10.65 80 ;
        RECT 9.375 78.15 9.875 80 ;
        RECT 8.6 78.15 9.1 80 ;
        RECT 7.825 78.15 8.325 80 ;
        RECT 7.05 78.15 7.55 80 ;
      LAYER C1 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IA ;
        RECT 7.35 77.975 10.35 80 ;
    END
  END VESD0_B
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 233.145 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 116.65125 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 493.90125 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 95.645 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 337.235 LAYER IA ;
    ANTENNAPARTIALMETALAREA 294.725 LAYER IB ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 10.276288 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 12.59712 LAYER YX ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER XA ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A2 ;
    ANTENNADIFFAREA 163.4 LAYER C5 ;
    ANTENNADIFFAREA 163.4 LAYER C4 ;
    ANTENNADIFFAREA 163.4 LAYER C6 ;
    ANTENNADIFFAREA 163.4 LAYER IA ;
    ANTENNADIFFAREA 163.4 LAYER IB ;
    ANTENNADIFFAREA 163.4 LAYER C3 ;
    PORT
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.875 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.875 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 2.35 21.75 57.65 25.35 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END PAD_B
  PIN VESD2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.0832 LAYER AY ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    PORT
      LAYER M1 ;
        RECT 38.35 78.15 38.85 80 ;
        RECT 37.575 78.15 38.075 80 ;
        RECT 36.8 78.15 37.3 80 ;
        RECT 36.025 78.15 36.525 80 ;
        RECT 35.25 78.15 35.75 80 ;
      LAYER M2 ;
        RECT 38.35 78.15 38.85 80 ;
        RECT 37.575 78.15 38.075 80 ;
        RECT 36.8 78.15 37.3 80 ;
        RECT 36.025 78.15 36.525 80 ;
        RECT 35.25 78.15 35.75 80 ;
      LAYER C1 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IA ;
        RECT 35.55 77.975 38.55 80 ;
    END
  END VESD2_B
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_ANAIO_V

MACRO RIIO_EG1D80V_CUTB2B_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTB2B_V 0 0 ;
  SIZE 16 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_r VSS_R!" ;
    PORT
      LAYER IB ;
        RECT 10 73.45 16 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 10 59.35 16 62.95 ;
    END
  END VSS_R
  PIN VSSIO_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_r VSSIO_R!" ;
    PORT
      LAYER IB ;
        RECT 10 54.65 16 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 10 45.25 16 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 10 40.55 16 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 10 26.45 16 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 10 17.05 16 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 10 3.67 16 6.55 ;
    END
  END VSSIO_R
  PIN VSSIO_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_l VSSIO_L!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 6 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 6 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 6 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 6 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 6 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 6 6.55 ;
    END
  END VSSIO_L
  PIN VSS_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_l VSS_L!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 6 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 6 62.95 ;
    END
  END VSS_L
  OBS
    LAYER CA ;
      RECT 0 0 16 80 ;
    LAYER M1 ;
      RECT 0 0 16 80 ;
    LAYER V1 ;
      RECT 0 0 16 80 ;
    LAYER M2 ;
      RECT 0 0 16 80 ;
    LAYER A1 ;
      RECT 0 0 16 80 ;
    LAYER C2 ;
      RECT 0 0 16 80 ;
    LAYER IA ;
      RECT 0 0 16 80 ;
    LAYER XA ;
      RECT 0 0 16 80 ;
    LAYER YX ;
      RECT 0 0 16 80 ;
    LAYER IB ;
      RECT 0 0 16 80 ;
    LAYER CB ;
      RECT 0 0 16 80 ;
    LAYER AY ;
      RECT 0 0 16 80 ;
    LAYER C1 ;
      RECT 0 0 16 80 ;
    LAYER C5 ;
      RECT 0 0 16 80 ;
    LAYER C4 ;
      RECT 0 0 16 80 ;
    LAYER C3 ;
      RECT 0 0 16 80 ;
    LAYER A5 ;
      RECT 0 0 16 80 ;
    LAYER A4 ;
      RECT 0 0 16 80 ;
    LAYER A3 ;
      RECT 0 0 16 80 ;
    LAYER A2 ;
      RECT 0 0 16 80 ;
    LAYER C6 ;
      RECT 0 0 16 80 ;
  END
END RIIO_EG1D80V_CUTB2B_V

MACRO RIIO_EG1D80V_CUTBIAS_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTBIAS_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 4 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 4 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 4 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 4 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 4 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 4 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 4 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 4 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 4 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 4 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 4 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 4 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 4 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 4 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 4 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTBIAS_V

MACRO RIIO_EG1D80V_CUTCOREB2B_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCOREB2B_V 0 0 ;
  SIZE 16 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 16 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 16 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 16 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 16 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 16 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 16 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 16 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 16 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 16 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 16 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 16 6.55 ;
    END
  END VSSIO
  PIN VSS_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_r VSS_R!" ;
    PORT
      LAYER IB ;
        RECT 8.875 73.45 16 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 8.875 59.35 16 62.95 ;
    END
  END VSS_R
  PIN VSS_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_l VSS_L!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 7.125 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 7.125 62.95 ;
    END
  END VSS_L
  OBS
    LAYER CA ;
      RECT 0 0 16 80 ;
    LAYER M1 ;
      RECT 0 0 16 80 ;
    LAYER V1 ;
      RECT 0 0 16 80 ;
    LAYER M2 ;
      RECT 0 0 16 80 ;
    LAYER A1 ;
      RECT 0 0 16 80 ;
    LAYER C2 ;
      RECT 0 0 16 80 ;
    LAYER IA ;
      RECT 0 0 16 80 ;
    LAYER XA ;
      RECT 0 0 16 80 ;
    LAYER YX ;
      RECT 0 0 16 80 ;
    LAYER IB ;
      RECT 0 0 16 80 ;
    LAYER CB ;
      RECT 0 0 16 80 ;
    LAYER AY ;
      RECT 0 0 16 80 ;
    LAYER C1 ;
      RECT 0 0 16 80 ;
    LAYER C5 ;
      RECT 0 0 16 80 ;
    LAYER C4 ;
      RECT 0 0 16 80 ;
    LAYER C3 ;
      RECT 0 0 16 80 ;
    LAYER A5 ;
      RECT 0 0 16 80 ;
    LAYER A4 ;
      RECT 0 0 16 80 ;
    LAYER A3 ;
      RECT 0 0 16 80 ;
    LAYER A2 ;
      RECT 0 0 16 80 ;
    LAYER C6 ;
      RECT 0 0 16 80 ;
  END
END RIIO_EG1D80V_CUTCOREB2B_V

MACRO RIIO_EG1D80V_CUTCOREPWR_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCOREPWR_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 4 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 4 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 4 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 4 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 4 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 4 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 4 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 4 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 4 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 4 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 4 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 4 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 4 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTCOREPWR_V

MACRO RIIO_EG1D80V_CUTCORE_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCORE_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 4 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 4 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 4 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 4 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 4 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 4 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 4 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 4 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 4 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 4 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 4 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTCORE_V

MACRO RIIO_EG1D80V_CUTIOB2B_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIOB2B_V 0 0 ;
  SIZE 16 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 16 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 16 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 16 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 16 67.65 ;
    END
  END VDD
  PIN VSSIO_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_l VSSIO_L!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 6 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 6 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 6 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 6 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 6 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 6 6.55 ;
    END
  END VSSIO_L
  PIN VSSIO_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_r VSSIO_R!" ;
    PORT
      LAYER IB ;
        RECT 10 54.65 16 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 10 45.25 16 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 10 40.55 16 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 10 26.45 16 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 10 17.05 16 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 10 3.67 16 6.55 ;
    END
  END VSSIO_R
  OBS
    LAYER CA ;
      RECT 0 0 16 80 ;
    LAYER M1 ;
      RECT 0 0 16 80 ;
    LAYER V1 ;
      RECT 0 0 16 80 ;
    LAYER M2 ;
      RECT 0 0 16 80 ;
    LAYER A1 ;
      RECT 0 0 16 80 ;
    LAYER C2 ;
      RECT 0 0 16 80 ;
    LAYER IA ;
      RECT 0 0 16 80 ;
    LAYER XA ;
      RECT 0 0 16 80 ;
    LAYER YX ;
      RECT 0 0 16 80 ;
    LAYER IB ;
      RECT 0 0 16 80 ;
    LAYER CB ;
      RECT 0 0 16 80 ;
    LAYER AY ;
      RECT 0 0 16 80 ;
    LAYER C1 ;
      RECT 0 0 16 80 ;
    LAYER C5 ;
      RECT 0 0 16 80 ;
    LAYER C4 ;
      RECT 0 0 16 80 ;
    LAYER C3 ;
      RECT 0 0 16 80 ;
    LAYER A5 ;
      RECT 0 0 16 80 ;
    LAYER A4 ;
      RECT 0 0 16 80 ;
    LAYER A3 ;
      RECT 0 0 16 80 ;
    LAYER A2 ;
      RECT 0 0 16 80 ;
    LAYER C6 ;
      RECT 0 0 16 80 ;
  END
END RIIO_EG1D80V_CUTIOB2B_V

MACRO RIIO_EG1D80V_CUTIOPWR_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIOPWR_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 4 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 4 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 4 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 4 67.65 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 4 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 4 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 4 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 4 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 4 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 4 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTIOPWR_V

MACRO RIIO_EG1D80V_CUTIO_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIO_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 4 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 4 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 4 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 4 67.65 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTIO_V

MACRO RIIO_EG1D80V_CUTPWR_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTPWR_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 4 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 4 62.95 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 4 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 4 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 4 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 4 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 4 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 4 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUTPWR_V

MACRO RIIO_EG1D80V_CUT_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUT_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_CUT_V

MACRO RIIO_EG1D80V_FILL16B2B_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL16B2B_V 0 0 ;
  SIZE 16 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 16 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 16 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 16 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 16 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 16 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 16 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 16 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 16 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 16 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 16 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 16 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 16 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 16 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 16 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 16 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 16 80 ;
    LAYER M1 ;
      RECT 0 0 16 80 ;
    LAYER V1 ;
      RECT 0 0 16 80 ;
    LAYER M2 ;
      RECT 0 0 16 80 ;
    LAYER A1 ;
      RECT 0 0 16 80 ;
    LAYER C2 ;
      RECT 0 0 16 80 ;
    LAYER IA ;
      RECT 0 0 16 80 ;
    LAYER XA ;
      RECT 0 0 16 80 ;
    LAYER YX ;
      RECT 0 0 16 80 ;
    LAYER IB ;
      RECT 0 0 16 80 ;
    LAYER CB ;
      RECT 0 0 16 80 ;
    LAYER AY ;
      RECT 0 0 16 80 ;
    LAYER C1 ;
      RECT 0 0 16 80 ;
    LAYER C5 ;
      RECT 0 0 16 80 ;
    LAYER C4 ;
      RECT 0 0 16 80 ;
    LAYER C3 ;
      RECT 0 0 16 80 ;
    LAYER A5 ;
      RECT 0 0 16 80 ;
    LAYER A4 ;
      RECT 0 0 16 80 ;
    LAYER A3 ;
      RECT 0 0 16 80 ;
    LAYER A2 ;
      RECT 0 0 16 80 ;
    LAYER C6 ;
      RECT 0 0 16 80 ;
  END
END RIIO_EG1D80V_FILL16B2B_V

MACRO RIIO_EG1D80V_FILL16_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL16_V 0 0 ;
  SIZE 16 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 16 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 16 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 16 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 16 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 16 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 16 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 16 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 16 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 16 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 16 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 16 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 16 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 16 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 16 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 16 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 16 80 ;
    LAYER M1 ;
      RECT 0 0 16 80 ;
    LAYER V1 ;
      RECT 0 0 16 80 ;
    LAYER M2 ;
      RECT 0 0 16 80 ;
    LAYER A1 ;
      RECT 0 0 16 80 ;
    LAYER C2 ;
      RECT 0 0 16 80 ;
    LAYER IA ;
      RECT 0 0 16 80 ;
    LAYER XA ;
      RECT 0 0 16 80 ;
    LAYER YX ;
      RECT 0 0 16 80 ;
    LAYER IB ;
      RECT 0 0 16 80 ;
    LAYER CB ;
      RECT 0 0 16 80 ;
    LAYER AY ;
      RECT 0 0 16 80 ;
    LAYER C1 ;
      RECT 0 0 16 80 ;
    LAYER C5 ;
      RECT 0 0 16 80 ;
    LAYER C4 ;
      RECT 0 0 16 80 ;
    LAYER C3 ;
      RECT 0 0 16 80 ;
    LAYER A5 ;
      RECT 0 0 16 80 ;
    LAYER A4 ;
      RECT 0 0 16 80 ;
    LAYER A3 ;
      RECT 0 0 16 80 ;
    LAYER A2 ;
      RECT 0 0 16 80 ;
    LAYER C6 ;
      RECT 0 0 16 80 ;
  END
END RIIO_EG1D80V_FILL16_V

MACRO RIIO_EG1D80V_FILL1_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL1_V 0 0 ;
  SIZE 1 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 1 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 1 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 1 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 1 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 1 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 1 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 1 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 1 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 1 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 1 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 1 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 1 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 1 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 1 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 1 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 1 80 ;
    LAYER M1 ;
      RECT 0 0 1 80 ;
    LAYER V1 ;
      RECT 0 0 1 80 ;
    LAYER M2 ;
      RECT 0 0 1 80 ;
    LAYER A1 ;
      RECT 0 0 1 80 ;
    LAYER C2 ;
      RECT 0 0 1 80 ;
    LAYER IA ;
      RECT 0 0 1 80 ;
    LAYER XA ;
      RECT 0 0 1 80 ;
    LAYER YX ;
      RECT 0 0 1 80 ;
    LAYER IB ;
      RECT 0 0 1 80 ;
    LAYER CB ;
      RECT 0 0 1 80 ;
    LAYER AY ;
      RECT 0 0 1 80 ;
    LAYER C1 ;
      RECT 0 0 1 80 ;
    LAYER C5 ;
      RECT 0 0 1 80 ;
    LAYER C4 ;
      RECT 0 0 1 80 ;
    LAYER C3 ;
      RECT 0 0 1 80 ;
    LAYER A5 ;
      RECT 0 0 1 80 ;
    LAYER A4 ;
      RECT 0 0 1 80 ;
    LAYER A3 ;
      RECT 0 0 1 80 ;
    LAYER A2 ;
      RECT 0 0 1 80 ;
    LAYER C6 ;
      RECT 0 0 1 80 ;
  END
END RIIO_EG1D80V_FILL1_V

MACRO RIIO_EG1D80V_FILL2_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL2_V 0 0 ;
  SIZE 2 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 2 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 2 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 2 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 2 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 2 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 2 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 2 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 2 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 2 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 2 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 2 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 2 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 2 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 2 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 2 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 2 80 ;
    LAYER M1 ;
      RECT 0 0 2 80 ;
    LAYER V1 ;
      RECT 0 0 2 80 ;
    LAYER M2 ;
      RECT 0 0 2 80 ;
    LAYER A1 ;
      RECT 0 0 2 80 ;
    LAYER C2 ;
      RECT 0 0 2 80 ;
    LAYER IA ;
      RECT 0 0 2 80 ;
    LAYER XA ;
      RECT 0 0 2 80 ;
    LAYER YX ;
      RECT 0 0 2 80 ;
    LAYER IB ;
      RECT 0 0 2 80 ;
    LAYER CB ;
      RECT 0 0 2 80 ;
    LAYER AY ;
      RECT 0 0 2 80 ;
    LAYER C1 ;
      RECT 0 0 2 80 ;
    LAYER C5 ;
      RECT 0 0 2 80 ;
    LAYER C4 ;
      RECT 0 0 2 80 ;
    LAYER C3 ;
      RECT 0 0 2 80 ;
    LAYER A5 ;
      RECT 0 0 2 80 ;
    LAYER A4 ;
      RECT 0 0 2 80 ;
    LAYER A3 ;
      RECT 0 0 2 80 ;
    LAYER A2 ;
      RECT 0 0 2 80 ;
    LAYER C6 ;
      RECT 0 0 2 80 ;
  END
END RIIO_EG1D80V_FILL2_V

MACRO RIIO_EG1D80V_FILL32_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL32_V 0 0 ;
  SIZE 32 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 32 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 32 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 32 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 32 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 32 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 32 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 32 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 32 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 32 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 32 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 32 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 32 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 32 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 32 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 32 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 32 80 ;
    LAYER M1 ;
      RECT 0 0 32 80 ;
    LAYER V1 ;
      RECT 0 0 32 80 ;
    LAYER M2 ;
      RECT 0 0 32 80 ;
    LAYER A1 ;
      RECT 0 0 32 80 ;
    LAYER C2 ;
      RECT 0 0 32 80 ;
    LAYER IA ;
      RECT 0 0 32 80 ;
    LAYER XA ;
      RECT 0 0 32 80 ;
    LAYER YX ;
      RECT 0 0 32 80 ;
    LAYER IB ;
      RECT 0 0 32 80 ;
    LAYER CB ;
      RECT 0 0 32 80 ;
    LAYER AY ;
      RECT 0 0 32 80 ;
    LAYER C1 ;
      RECT 0 0 32 80 ;
    LAYER C5 ;
      RECT 0 0 32 80 ;
    LAYER C4 ;
      RECT 0 0 32 80 ;
    LAYER C3 ;
      RECT 0 0 32 80 ;
    LAYER A5 ;
      RECT 0 0 32 80 ;
    LAYER A4 ;
      RECT 0 0 32 80 ;
    LAYER A3 ;
      RECT 0 0 32 80 ;
    LAYER A2 ;
      RECT 0 0 32 80 ;
    LAYER C6 ;
      RECT 0 0 32 80 ;
  END
END RIIO_EG1D80V_FILL32_V

MACRO RIIO_EG1D80V_FILL4_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL4_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 4 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 4 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 4 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 4 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 4 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 4 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 4 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 4 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 4 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 4 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 4 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 4 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 4 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 4 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 4 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_FILL4_V

MACRO RIIO_EG1D80V_FILL8_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL8_V 0 0 ;
  SIZE 8 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 8 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 8 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 8 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 8 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 8 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 8 6.55 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 8 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 8 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 8 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 8 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 8 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 8 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 8 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 8 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 8 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 8 80 ;
    LAYER M1 ;
      RECT 0 0 8 80 ;
    LAYER V1 ;
      RECT 0 0 8 80 ;
    LAYER M2 ;
      RECT 0 0 8 80 ;
    LAYER A1 ;
      RECT 0 0 8 80 ;
    LAYER C2 ;
      RECT 0 0 8 80 ;
    LAYER IA ;
      RECT 0 0 8 80 ;
    LAYER XA ;
      RECT 0 0 8 80 ;
    LAYER YX ;
      RECT 0 0 8 80 ;
    LAYER IB ;
      RECT 0 0 8 80 ;
    LAYER CB ;
      RECT 0 0 8 80 ;
    LAYER AY ;
      RECT 0 0 8 80 ;
    LAYER C1 ;
      RECT 0 0 8 80 ;
    LAYER C5 ;
      RECT 0 0 8 80 ;
    LAYER C4 ;
      RECT 0 0 8 80 ;
    LAYER C3 ;
      RECT 0 0 8 80 ;
    LAYER A5 ;
      RECT 0 0 8 80 ;
    LAYER A4 ;
      RECT 0 0 8 80 ;
    LAYER A3 ;
      RECT 0 0 8 80 ;
    LAYER A2 ;
      RECT 0 0 8 80 ;
    LAYER C6 ;
      RECT 0 0 8 80 ;
  END
END RIIO_EG1D80V_FILL8_V

MACRO RIIO_EG1D80V_POR_IO_V1D0_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_POR_IO_V1D0_V 0 0 ;
  SIZE 8 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER C2 ;
        RECT 0 37.075 8 39.575 ;
    END
    PORT
      LAYER IB ;
        RECT 0 54.65 8 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 8 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 8 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 8 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 8 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 8 6.55 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 8 77.05 ;
      LAYER C2 ;
        RECT 0 74.575 8 77.075 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 8 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 8 72.35 ;
      LAYER C2 ;
        RECT 0 70.825 8 73.325 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 8 67.65 ;
    END
  END VDD
  PIN VDDIO_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio_por VDDIO_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 1.25 33.325 1.75 80 ;
    END
  END VDDIO_POR
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 8 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 8 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 8 34.75 ;
      LAYER C2 ;
        RECT 0 33.325 8 35.825 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 8 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 8 11.25 ;
    END
  END VDDIO
  PIN VSSIO_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_por VSSIO_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 2.25 33.325 2.75 80 ;
    END
  END VSSIO_POR
  PIN POR_N_CORE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.5875 LAYER C1 ;
    ANTENNADIFFAREA 0.3135 LAYER C1 ;
    PORT
      LAYER C1 ;
        RECT 6.25 79.5 6.75 80 ;
    END
  END POR_N_CORE_O
  PIN VDD_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd_por VDD_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 5.25 70.825 5.75 80 ;
    END
  END VDD_POR
  PIN VSS_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_por VSS_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C1 ;
        RECT 4.25 70.825 4.75 80 ;
    END
  END VSS_POR
  OBS
    LAYER CA ;
      RECT 0 0 8 80 ;
    LAYER M1 ;
      RECT 0 0 8 80 ;
    LAYER V1 ;
      RECT 0 0 8 80 ;
    LAYER M2 ;
      RECT 0 0 8 80 ;
    LAYER A1 ;
      RECT 0 0 8 80 ;
    LAYER C2 ;
      RECT 0 0 8 80 ;
    LAYER IA ;
      RECT 0 0 8 80 ;
    LAYER XA ;
      RECT 0 0 8 80 ;
    LAYER YX ;
      RECT 0 0 8 80 ;
    LAYER IB ;
      RECT 0 0 8 80 ;
    LAYER CB ;
      RECT 0 0 8 80 ;
    LAYER AY ;
      RECT 0 0 8 80 ;
    LAYER C1 ;
      RECT 0 0 8 80 ;
    LAYER C5 ;
      RECT 0 0 8 80 ;
    LAYER C4 ;
      RECT 0 0 8 80 ;
    LAYER C3 ;
      RECT 0 0 8 80 ;
    LAYER A5 ;
      RECT 0 0 8 80 ;
    LAYER A4 ;
      RECT 0 0 8 80 ;
    LAYER A3 ;
      RECT 0 0 8 80 ;
    LAYER A2 ;
      RECT 0 0 8 80 ;
    LAYER C6 ;
      RECT 0 0 8 80 ;
  END
END RIIO_EG1D80V_POR_IO_V1D0_V

MACRO RIIO_EG1D80V_RAILSHORT_GND_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_GND_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 4 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 4 62.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 54.65 4 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 4 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 4 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 4 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 4 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 4 6.55 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 4 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 4 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 4 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 4 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 4 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 4 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 4 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_RAILSHORT_GND_V

MACRO RIIO_EG1D80V_RAILSHORT_PG_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_PG_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 4 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 4 62.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 54.65 4 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 4 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 4 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 4 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 4 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 4 6.55 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 4 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 4 67.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.95 4 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 4 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 4 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 4 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 4 11.25 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_RAILSHORT_PG_V

MACRO RIIO_EG1D80V_RAILSHORT_PWR_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_PWR_V 0 0 ;
  SIZE 4 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 4 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 4 67.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.95 4 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 4 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 4 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 4 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 4 11.25 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 4 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 4 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 4 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 4 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 4 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 4 6.55 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 4 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 4 62.95 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 4 80 ;
    LAYER M1 ;
      RECT 0 0 4 80 ;
    LAYER V1 ;
      RECT 0 0 4 80 ;
    LAYER M2 ;
      RECT 0 0 4 80 ;
    LAYER A1 ;
      RECT 0 0 4 80 ;
    LAYER C2 ;
      RECT 0 0 4 80 ;
    LAYER IA ;
      RECT 0 0 4 80 ;
    LAYER XA ;
      RECT 0 0 4 80 ;
    LAYER YX ;
      RECT 0 0 4 80 ;
    LAYER IB ;
      RECT 0 0 4 80 ;
    LAYER CB ;
      RECT 0 0 4 80 ;
    LAYER AY ;
      RECT 0 0 4 80 ;
    LAYER C1 ;
      RECT 0 0 4 80 ;
    LAYER C5 ;
      RECT 0 0 4 80 ;
    LAYER C4 ;
      RECT 0 0 4 80 ;
    LAYER C3 ;
      RECT 0 0 4 80 ;
    LAYER A5 ;
      RECT 0 0 4 80 ;
    LAYER A4 ;
      RECT 0 0 4 80 ;
    LAYER A3 ;
      RECT 0 0 4 80 ;
    LAYER A2 ;
      RECT 0 0 4 80 ;
    LAYER C6 ;
      RECT 0 0 4 80 ;
  END
END RIIO_EG1D80V_RAILSHORT_PWR_V

MACRO RIIO_EG1D80V_VDD04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
    END
    PORT
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
    END
    PORT
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
    END
    PORT
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
    END
    PORT
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
    END
    PORT
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDD04_V

MACRO RIIO_EG1D80V_VDDIOX_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDIOX_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSSIOX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssiox VSSIOX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C2 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C1 ;
        RECT 9.837 79.19 12.662 80 ;
      LAYER M2 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER M1 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C2 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C1 ;
        RECT 47.337 79.19 50.162 80 ;
      LAYER M2 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER M1 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
  END VSSIOX
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDDIOX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddiox VDDIOX!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VDDIOX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDIOX_V

MACRO RIIO_EG1D80V_VDDIO_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDIO_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDIO_V

MACRO RIIO_EG1D80V_VDDQ04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VDDQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDQ04_V

MACRO RIIO_EG1D80V_VDDQ_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VDDQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDQ_HVT_V

MACRO RIIO_EG1D80V_VDDQ_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VDDQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDQ_RVT_V

MACRO RIIO_EG1D80V_VDDX04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C2 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C1 ;
        RECT 9.837 79.19 12.662 80 ;
      LAYER M2 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER M1 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C2 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C1 ;
        RECT 47.337 79.19 50.162 80 ;
      LAYER M2 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER M1 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDX04_V

MACRO RIIO_EG1D80V_VDDX_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C2 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C1 ;
        RECT 9.837 79.19 12.662 80 ;
      LAYER M2 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER M1 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C2 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C1 ;
        RECT 47.337 79.19 50.162 80 ;
      LAYER M2 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER M1 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDX_HVT_V

MACRO RIIO_EG1D80V_VDDX_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C2 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C1 ;
        RECT 9.837 79.19 12.662 80 ;
      LAYER M2 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER M1 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C2 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C1 ;
        RECT 47.337 79.19 50.162 80 ;
      LAYER M2 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER M1 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDDX_RVT_V

MACRO RIIO_EG1D80V_VDD_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDD_HVT_V

MACRO RIIO_EG1D80V_VDD_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VDD_RVT_V

MACRO RIIO_EG1D80V_VNWINT_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNWINT_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VNWINT_HVT_V

MACRO RIIO_EG1D80V_VNWINT_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNWINT_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VNWINT_RVT_V

MACRO RIIO_EG1D80V_VNW_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNW_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VNW_V

MACRO RIIO_EG1D80V_VPWINT_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPWINT_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VPWINT_HVT_V

MACRO RIIO_EG1D80V_VPWINT_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPWINT_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VPWINT_RVT_V

MACRO RIIO_EG1D80V_VPW_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPW_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VPW_V

MACRO RIIO_EG1D80V_VSS04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
    END
    PORT
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
    END
    PORT
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
    END
    PORT
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
    END
    PORT
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
    END
    PORT
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSS04_V

MACRO RIIO_EG1D80V_VSSIOX_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSIOX_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSIOX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssiox VSSIOX!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C2 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C1 ;
        RECT 9.837 79.19 12.662 80 ;
      LAYER M2 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER M1 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C2 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C1 ;
        RECT 47.337 79.19 50.162 80 ;
      LAYER M2 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER M1 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSSIOX
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDDIOX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddiox VDDIOX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
  END VDDIOX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSIOX_V

MACRO RIIO_EG1D80V_VSSIO_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSIO_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSIO_V

MACRO RIIO_EG1D80V_VSSQ04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDQ
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSSQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSQ04_V

MACRO RIIO_EG1D80V_VSSQ_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSSQ
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSQ_HVT_V

MACRO RIIO_EG1D80V_VSSQ_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSSQ
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDQ
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSQ_RVT_V

MACRO RIIO_EG1D80V_VSSX04_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX04_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C2 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C1 ;
        RECT 9.837 79.19 12.662 80 ;
      LAYER M2 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER M1 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C2 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C1 ;
        RECT 47.337 79.19 50.162 80 ;
      LAYER M2 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER M1 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSX04_V

MACRO RIIO_EG1D80V_VSSX_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C2 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C1 ;
        RECT 9.837 79.19 12.662 80 ;
      LAYER M2 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER M1 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C2 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C1 ;
        RECT 47.337 79.19 50.162 80 ;
      LAYER M2 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER M1 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSX_HVT_V

MACRO RIIO_EG1D80V_VSSX_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C2 ;
        RECT 17.5 78.15 20 80 ;
      LAYER C1 ;
        RECT 17.337 79.19 20.162 80 ;
      LAYER M2 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
      LAYER M1 ;
        RECT 19.662 79.19 20.162 80 ;
        RECT 18.887 79.19 19.387 80 ;
        RECT 18.112 79.19 18.612 80 ;
        RECT 17.337 79.19 17.837 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C2 ;
        RECT 40 78.15 42.5 80 ;
      LAYER C1 ;
        RECT 39.837 79.19 42.662 80 ;
      LAYER M2 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
      LAYER M1 ;
        RECT 42.162 79.19 42.662 80 ;
        RECT 41.387 79.19 41.887 80 ;
        RECT 40.612 79.19 41.112 80 ;
        RECT 39.837 79.19 40.337 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C2 ;
        RECT 10 78.15 12.5 80 ;
      LAYER C1 ;
        RECT 9.837 79.19 12.662 80 ;
      LAYER M2 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER M1 ;
        RECT 12.162 79.19 12.662 80 ;
        RECT 11.387 79.19 11.887 80 ;
        RECT 10.612 79.19 11.112 80 ;
        RECT 9.837 79.19 10.337 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C2 ;
        RECT 25 78.15 27.5 80 ;
      LAYER C1 ;
        RECT 24.837 79.19 27.662 80 ;
      LAYER M2 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER M1 ;
        RECT 27.162 79.19 27.662 80 ;
        RECT 26.387 79.19 26.887 80 ;
        RECT 25.612 79.19 26.112 80 ;
        RECT 24.837 79.19 25.337 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C2 ;
        RECT 32.5 78.15 35 80 ;
      LAYER C1 ;
        RECT 32.337 79.19 35.162 80 ;
      LAYER M2 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER M1 ;
        RECT 34.662 79.19 35.162 80 ;
        RECT 33.887 79.19 34.387 80 ;
        RECT 33.112 79.19 33.612 80 ;
        RECT 32.337 79.19 32.837 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C2 ;
        RECT 47.5 78.15 50 80 ;
      LAYER C1 ;
        RECT 47.337 79.19 50.162 80 ;
      LAYER M2 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER M1 ;
        RECT 49.662 79.19 50.162 80 ;
        RECT 48.887 79.19 49.387 80 ;
        RECT 48.112 79.19 48.612 80 ;
        RECT 47.337 79.19 47.837 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C2 ;
        RECT 21.25 78.15 23.75 80 ;
      LAYER C1 ;
        RECT 21.087 79.19 23.912 80 ;
      LAYER M2 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
      LAYER M1 ;
        RECT 23.412 79.19 23.912 80 ;
        RECT 22.637 79.19 23.137 80 ;
        RECT 21.862 79.19 22.362 80 ;
        RECT 21.087 79.19 21.587 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C2 ;
        RECT 28.75 78.15 31.25 80 ;
      LAYER C1 ;
        RECT 28.587 79.19 31.412 80 ;
      LAYER M2 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
      LAYER M1 ;
        RECT 30.912 79.19 31.412 80 ;
        RECT 30.137 79.19 30.637 80 ;
        RECT 29.362 79.19 29.862 80 ;
        RECT 28.587 79.19 29.087 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C2 ;
        RECT 36.25 78.15 38.75 80 ;
      LAYER C1 ;
        RECT 36.087 79.19 38.912 80 ;
      LAYER M2 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
      LAYER M1 ;
        RECT 38.412 79.19 38.912 80 ;
        RECT 37.637 79.19 38.137 80 ;
        RECT 36.862 79.19 37.362 80 ;
        RECT 36.087 79.19 36.587 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C2 ;
        RECT 13.75 78.15 16.25 80 ;
      LAYER C1 ;
        RECT 13.587 79.19 16.412 80 ;
      LAYER M2 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER M1 ;
        RECT 15.912 79.19 16.412 80 ;
        RECT 15.137 79.19 15.637 80 ;
        RECT 14.362 79.19 14.862 80 ;
        RECT 13.587 79.19 14.087 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C2 ;
        RECT 43.75 78.15 46.25 80 ;
      LAYER C1 ;
        RECT 43.587 79.19 46.412 80 ;
      LAYER M2 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER M1 ;
        RECT 45.912 79.19 46.412 80 ;
        RECT 45.137 79.19 45.637 80 ;
        RECT 44.362 79.19 44.862 80 ;
        RECT 43.587 79.19 44.087 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSSX_RVT_V

MACRO RIIO_EG1D80V_VSS_HVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS_HVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSS_HVT_V

MACRO RIIO_EG1D80V_VSS_RVT_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS_RVT_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
    END
    PORT
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
    END
    PORT
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
    END
    PORT
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
    END
    PORT
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
    END
    PORT
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
    END
    PORT
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
    END
    PORT
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
    END
    PORT
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
    END
    PORT
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
    END
    PORT
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSS_RVT_V

MACRO RIIO_EG1D80V_VSUP_CORE_GND_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_GND_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
    END
    PORT
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
    END
    PORT
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
    END
    PORT
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
    END
    PORT
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
    END
    PORT
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSUP
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_CORE_GND_V

MACRO RIIO_EG1D80V_VSUP_CORE_PWR_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_PWR_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
    END
    PORT
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
    END
    PORT
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
    END
    PORT
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
    END
    PORT
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
    END
    PORT
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSUP
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_CORE_PWR_V

MACRO RIIO_EG1D80V_VSUP_CORE_SIG_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_SIG_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1201.173 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 4.4055 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 514.88 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 1152.81 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 610.4525 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 944.67 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 770.45 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1268.18 LAYER IA ;
    ANTENNAPARTIALMETALAREA 398.14 LAYER IB ;
    ANTENNAPARTIALMETALAREA 4.554 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 18.283584 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 1.792 LAYER AY ;
    ANTENNAPARTIALCUTAREA 16.239168 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 26.515456 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 62.9856 LAYER YX ;
    ANTENNAPARTIALCUTAREA 40.310784 LAYER XA ;
    ANTENNAPARTIALCUTAREA 1.92 LAYER V1 ;
    ANTENNADIFFAREA 150.1 LAYER C3 ;
    ANTENNADIFFAREA 150.1 LAYER C2 ;
    ANTENNADIFFAREA 150.1 LAYER C4 ;
    ANTENNADIFFAREA 150.1 LAYER C5 ;
    ANTENNADIFFAREA 150.1 LAYER C6 ;
    ANTENNADIFFAREA 150.1 LAYER IA ;
    ANTENNADIFFAREA 150.1 LAYER IB ;
    ANTENNADIFFAREA 150.1 LAYER C1 ;
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
        RECT 2.65 79.19 5.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 2.35 21.75 57.65 25.35 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END VSUP
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_CORE_SIG_V

MACRO RIIO_EG1D80V_VSUP_IO_GND_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_GND_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
    END
    PORT
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
    END
    PORT
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
    END
    PORT
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
    END
    PORT
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
    END
    PORT
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSUP
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_IO_GND_V

MACRO RIIO_EG1D80V_VSUP_IO_PWR_V
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_PWR_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IA ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C2 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C1 ;
        RECT 2.65 79.19 5.65 80 ;
      LAYER M2 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER M1 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 2.35 0 5.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER IA ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C6 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C5 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C4 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C3 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C2 ;
        RECT 7.35 78.15 10.35 80 ;
      LAYER C1 ;
        RECT 7.35 79.19 10.35 80 ;
      LAYER M2 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
      LAYER M1 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER IA ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C6 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C5 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C4 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C3 ;
        RECT 7.05 0 10.65 1.85 ;
      LAYER C2 ;
        RECT 7.05 0 10.65 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER IA ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C6 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C5 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C4 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C3 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C2 ;
        RECT 12.05 78.15 15.05 80 ;
      LAYER C1 ;
        RECT 12.05 79.19 15.05 80 ;
      LAYER M2 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
      LAYER M1 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
    END
    PORT
      LAYER IB ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER IA ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C6 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C5 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C4 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C3 ;
        RECT 11.75 0 15.35 1.85 ;
      LAYER C2 ;
        RECT 11.75 0 15.35 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER IA ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C6 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C5 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C4 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C3 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C2 ;
        RECT 16.75 78.15 19.75 80 ;
      LAYER C1 ;
        RECT 16.75 79.19 19.75 80 ;
      LAYER M2 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
      LAYER M1 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
    END
    PORT
      LAYER IB ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER IA ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C6 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C5 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C4 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C3 ;
        RECT 16.45 0 20.05 1.85 ;
      LAYER C2 ;
        RECT 16.45 0 20.05 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER IA ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C6 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C5 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C4 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C3 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C2 ;
        RECT 21.45 78.15 24.45 80 ;
      LAYER C1 ;
        RECT 21.45 79.19 24.45 80 ;
      LAYER M2 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
      LAYER M1 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER IA ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C6 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C5 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C4 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C3 ;
        RECT 21.15 0 24.75 1.85 ;
      LAYER C2 ;
        RECT 21.15 0 24.75 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER IA ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C6 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C5 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C4 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C3 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C2 ;
        RECT 26.15 78.15 29.15 80 ;
      LAYER C1 ;
        RECT 26.15 79.19 29.15 80 ;
      LAYER M2 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
      LAYER M1 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
    END
    PORT
      LAYER IB ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER IA ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C6 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C5 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C4 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C3 ;
        RECT 25.85 0 29.45 1.85 ;
      LAYER C2 ;
        RECT 25.85 0 29.45 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER IA ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C6 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C5 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C4 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C3 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C2 ;
        RECT 30.85 78.15 33.85 80 ;
      LAYER C1 ;
        RECT 30.85 79.19 33.85 80 ;
      LAYER M2 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
      LAYER M1 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
    END
    PORT
      LAYER IB ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER IA ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C6 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C5 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C4 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C3 ;
        RECT 30.55 0 34.15 1.85 ;
      LAYER C2 ;
        RECT 30.55 0 34.15 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER IA ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C6 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C5 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C4 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C3 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C2 ;
        RECT 35.55 78.15 38.55 80 ;
      LAYER C1 ;
        RECT 35.55 79.19 38.55 80 ;
      LAYER M2 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
      LAYER M1 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
    END
    PORT
      LAYER IB ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER IA ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C6 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C5 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C4 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C3 ;
        RECT 35.25 0 38.85 1.85 ;
      LAYER C2 ;
        RECT 35.25 0 38.85 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER IA ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C6 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C5 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C4 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C3 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C2 ;
        RECT 40.25 78.15 43.25 80 ;
      LAYER C1 ;
        RECT 40.25 79.19 43.25 80 ;
      LAYER M2 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
      LAYER M1 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
    END
    PORT
      LAYER IB ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER IA ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C6 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C5 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C4 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C3 ;
        RECT 39.95 0 43.55 1.85 ;
      LAYER C2 ;
        RECT 39.95 0 43.55 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER IA ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C6 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C5 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C4 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C3 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C2 ;
        RECT 44.95 78.15 47.95 80 ;
      LAYER C1 ;
        RECT 44.95 79.19 47.95 80 ;
      LAYER M2 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
      LAYER M1 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
    END
    PORT
      LAYER IB ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER IA ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C6 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C5 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C4 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C3 ;
        RECT 44.65 0 48.25 1.85 ;
      LAYER C2 ;
        RECT 44.65 0 48.25 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER IA ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C6 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C5 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C4 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C3 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C2 ;
        RECT 49.65 78.15 52.65 80 ;
      LAYER C1 ;
        RECT 49.65 79.19 52.65 80 ;
      LAYER M2 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
      LAYER M1 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
    END
    PORT
      LAYER IB ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER IA ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C6 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C5 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C4 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C3 ;
        RECT 49.35 0 52.95 1.85 ;
      LAYER C2 ;
        RECT 49.35 0 52.95 1.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
    END
    PORT
      LAYER IB ;
        RECT 2.35 21.75 57.65 25.35 ;
    END
    PORT
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
    END
  END VSUP
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_IO_PWR_V

MACRO RIIO_EG1D80V_VSUP_IO_SIG_V
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_SIG_V 0 0 ;
  SIZE 60 BY 80 ;
  SYMMETRY X Y ;
  SITE IO_NS_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1543.173 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 4.4055 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 654.255 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 1152.81 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 610.4525 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 944.67 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 770.45 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1268.18 LAYER IA ;
    ANTENNAPARTIALMETALAREA 397.03 LAYER IB ;
    ANTENNAPARTIALMETALAREA 4.554 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 23.58048 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 1.792 LAYER AY ;
    ANTENNAPARTIALCUTAREA 19.220608 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 26.515456 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 62.9856 LAYER YX ;
    ANTENNAPARTIALCUTAREA 40.310784 LAYER XA ;
    ANTENNAPARTIALCUTAREA 1.92 LAYER V1 ;
    ANTENNADIFFAREA 163.4 LAYER C3 ;
    ANTENNADIFFAREA 163.4 LAYER C2 ;
    ANTENNADIFFAREA 163.4 LAYER C4 ;
    ANTENNADIFFAREA 163.4 LAYER C5 ;
    ANTENNADIFFAREA 163.4 LAYER C6 ;
    ANTENNADIFFAREA 163.4 LAYER IA ;
    ANTENNADIFFAREA 163.4 LAYER IB ;
    ANTENNADIFFAREA 163.4 LAYER C1 ;
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER IA ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C6 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C5 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C4 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER C3 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER M1 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER C2 ;
        RECT 54.35 78.15 57.35 80 ;
        RECT 49.65 78.15 52.65 80 ;
        RECT 44.95 78.15 47.95 80 ;
        RECT 40.25 78.15 43.25 80 ;
        RECT 35.55 78.15 38.55 80 ;
        RECT 30.85 78.15 33.85 80 ;
        RECT 26.15 78.15 29.15 80 ;
        RECT 21.45 78.15 24.45 80 ;
        RECT 16.75 78.15 19.75 80 ;
        RECT 12.05 78.15 15.05 80 ;
        RECT 7.35 78.15 10.35 80 ;
        RECT 2.65 78.15 5.65 80 ;
      LAYER M2 ;
        RECT 57.15 79.19 57.65 80 ;
        RECT 56.375 79.19 56.875 80 ;
        RECT 55.6 79.19 56.1 80 ;
        RECT 54.825 79.19 55.325 80 ;
        RECT 54.05 79.19 54.55 80 ;
        RECT 52.45 79.19 52.95 80 ;
        RECT 51.675 79.19 52.175 80 ;
        RECT 50.9 79.19 51.4 80 ;
        RECT 50.125 79.19 50.625 80 ;
        RECT 49.35 79.19 49.85 80 ;
        RECT 47.75 79.19 48.25 80 ;
        RECT 46.975 79.19 47.475 80 ;
        RECT 46.2 79.19 46.7 80 ;
        RECT 45.425 79.19 45.925 80 ;
        RECT 44.65 79.19 45.15 80 ;
        RECT 43.05 79.19 43.55 80 ;
        RECT 42.275 79.19 42.775 80 ;
        RECT 41.5 79.19 42 80 ;
        RECT 40.725 79.19 41.225 80 ;
        RECT 39.95 79.19 40.45 80 ;
        RECT 38.35 79.19 38.85 80 ;
        RECT 37.575 79.19 38.075 80 ;
        RECT 36.8 79.19 37.3 80 ;
        RECT 36.025 79.19 36.525 80 ;
        RECT 35.25 79.19 35.75 80 ;
        RECT 33.65 79.19 34.15 80 ;
        RECT 32.875 79.19 33.375 80 ;
        RECT 32.1 79.19 32.6 80 ;
        RECT 31.325 79.19 31.825 80 ;
        RECT 30.55 79.19 31.05 80 ;
        RECT 28.95 79.19 29.45 80 ;
        RECT 28.175 79.19 28.675 80 ;
        RECT 27.4 79.19 27.9 80 ;
        RECT 26.625 79.19 27.125 80 ;
        RECT 25.85 79.19 26.35 80 ;
        RECT 24.25 79.19 24.75 80 ;
        RECT 23.475 79.19 23.975 80 ;
        RECT 22.7 79.19 23.2 80 ;
        RECT 21.925 79.19 22.425 80 ;
        RECT 21.15 79.19 21.65 80 ;
        RECT 19.55 79.19 20.05 80 ;
        RECT 18.775 79.19 19.275 80 ;
        RECT 18 79.19 18.5 80 ;
        RECT 17.225 79.19 17.725 80 ;
        RECT 16.45 79.19 16.95 80 ;
        RECT 14.85 79.19 15.35 80 ;
        RECT 14.075 79.19 14.575 80 ;
        RECT 13.3 79.19 13.8 80 ;
        RECT 12.525 79.19 13.025 80 ;
        RECT 11.75 79.19 12.25 80 ;
        RECT 10.15 79.19 10.65 80 ;
        RECT 9.375 79.19 9.875 80 ;
        RECT 8.6 79.19 9.1 80 ;
        RECT 7.825 79.19 8.325 80 ;
        RECT 7.05 79.19 7.55 80 ;
        RECT 5.45 79.19 5.95 80 ;
        RECT 4.675 79.19 5.175 80 ;
        RECT 3.9 79.19 4.4 80 ;
        RECT 3.125 79.19 3.625 80 ;
        RECT 2.35 79.19 2.85 80 ;
      LAYER C1 ;
        RECT 54.35 79.19 57.35 80 ;
        RECT 49.65 79.19 52.65 80 ;
        RECT 44.95 79.19 47.95 80 ;
        RECT 40.25 79.19 43.25 80 ;
        RECT 35.55 79.19 38.55 80 ;
        RECT 30.85 79.19 33.85 80 ;
        RECT 26.15 79.19 29.15 80 ;
        RECT 21.45 79.19 24.45 80 ;
        RECT 16.75 79.19 19.75 80 ;
        RECT 12.05 79.19 15.05 80 ;
        RECT 7.35 79.19 10.35 80 ;
        RECT 2.65 79.19 5.65 80 ;
    END
    PORT
      LAYER IB ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 2.35 21.75 57.65 25.35 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER IA ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C6 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C5 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C4 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C3 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
      LAYER C2 ;
        RECT 54.05 0 57.65 1.85 ;
        RECT 49.35 0 52.95 1.85 ;
        RECT 44.65 0 48.25 1.85 ;
        RECT 39.95 0 43.55 1.85 ;
        RECT 35.25 0 38.85 1.85 ;
        RECT 30.55 0 34.15 1.85 ;
        RECT 25.85 0 29.45 1.85 ;
        RECT 21.15 0 24.75 1.85 ;
        RECT 16.45 0 20.05 1.85 ;
        RECT 11.75 0 15.35 1.85 ;
        RECT 7.05 0 10.65 1.85 ;
        RECT 2.35 0 5.95 1.85 ;
    END
  END VSUP
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 0 54.65 60 58.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 45.25 60 48.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 40.55 60 44.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 26.45 60 30.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 17.05 60 20.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 3.67 60 6.55 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 0 68.75 60 72.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 64.05 60 67.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 0 73.45 60 77.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 59.35 60 62.95 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 0 49.95 60 53.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.85 60 39.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 31.15 60 34.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 12.35 60 15.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.65 60 11.25 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 60 80 ;
    LAYER M1 ;
      RECT 0 0 60 80 ;
    LAYER V1 ;
      RECT 0 0 60 80 ;
    LAYER M2 ;
      RECT 0 0 60 80 ;
    LAYER A1 ;
      RECT 0 0 60 80 ;
    LAYER C2 ;
      RECT 0 0 60 80 ;
    LAYER IA ;
      RECT 0 0 60 80 ;
    LAYER XA ;
      RECT 0 0 60 80 ;
    LAYER YX ;
      RECT 0 0 60 80 ;
    LAYER IB ;
      RECT 0 0 60 80 ;
    LAYER CB ;
      RECT 0 0 60 80 ;
    LAYER AY ;
      RECT 0 0 60 80 ;
    LAYER C1 ;
      RECT 0 0 60 80 ;
    LAYER C5 ;
      RECT 0 0 60 80 ;
    LAYER C4 ;
      RECT 0 0 60 80 ;
    LAYER C3 ;
      RECT 0 0 60 80 ;
    LAYER A5 ;
      RECT 0 0 60 80 ;
    LAYER A4 ;
      RECT 0 0 60 80 ;
    LAYER A3 ;
      RECT 0 0 60 80 ;
    LAYER A2 ;
      RECT 0 0 60 80 ;
    LAYER C6 ;
      RECT 0 0 60 80 ;
  END
END RIIO_EG1D80V_VSUP_IO_SIG_V

MACRO RIIO_EG1D80V_ANACORE_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ANACORE_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 95.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 567.2075 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 603.245 LAYER IA ;
    ANTENNAPARTIALMETALAREA 294.725 LAYER IB ;
    ANTENNAPARTIALMETALAREA 188.175 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 12.04192 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 11.54736 LAYER YX ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER XA ;
    ANTENNAPARTIALCUTAREA 4.232096 LAYER A2 ;
    ANTENNADIFFAREA 133.0532 LAYER C4 ;
    ANTENNADIFFAREA 133.0532 LAYER C3 ;
    ANTENNADIFFAREA 133.0532 LAYER C5 ;
    ANTENNADIFFAREA 133.0532 LAYER C6 ;
    ANTENNADIFFAREA 133.0532 LAYER IA ;
    ANTENNADIFFAREA 133.0532 LAYER IB ;
    ANTENNADIFFAREA 133.0532 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN VRES3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.735 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 79.654 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 93.78 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.4675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.3648 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 11.75 80 12.25 ;
        RECT 78.15 12.525 80 13.025 ;
        RECT 78.15 13.3 80 13.8 ;
        RECT 78.15 14.075 80 14.575 ;
        RECT 78.15 14.85 80 15.35 ;
      LAYER M2 ;
        RECT 78.15 11.75 80 12.25 ;
        RECT 78.15 12.525 80 13.025 ;
        RECT 78.15 13.3 80 13.8 ;
        RECT 78.15 14.075 80 14.575 ;
        RECT 78.15 14.85 80 15.35 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 77.975 12.05 80 15.05 ;
    END
  END VRES3_B
  PIN VESD0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 24.7745 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 93.505 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 49.35 80 49.85 ;
        RECT 78.15 50.125 80 50.625 ;
        RECT 78.15 50.9 80 51.4 ;
        RECT 78.15 51.675 80 52.175 ;
        RECT 78.15 52.45 80 52.95 ;
      LAYER M2 ;
        RECT 78.15 49.35 80 49.85 ;
        RECT 78.15 50.125 80 50.625 ;
        RECT 78.15 50.9 80 51.4 ;
        RECT 78.15 51.675 80 52.175 ;
        RECT 78.15 52.45 80 52.95 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 77.975 49.65 80 52.65 ;
    END
  END VESD0_B
  PIN VRES0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.235 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 36.0415 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 91.905 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.4675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.099 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.747296 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.6144 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.1664 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 44.65 80 45.15 ;
        RECT 78.15 45.425 80 45.925 ;
        RECT 78.15 46.2 80 46.7 ;
        RECT 78.15 46.975 80 47.475 ;
        RECT 78.15 47.75 80 48.25 ;
      LAYER M2 ;
        RECT 78.15 44.65 80 45.15 ;
        RECT 78.15 45.425 80 45.925 ;
        RECT 78.15 46.2 80 46.7 ;
        RECT 78.15 46.975 80 47.475 ;
        RECT 78.15 47.75 80 48.25 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 77.975 44.95 80 47.95 ;
    END
  END VRES0_B
  PIN VRES1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.235 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 22.887 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 87.235 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 39.95 80 40.45 ;
        RECT 78.15 40.725 80 41.225 ;
        RECT 78.15 41.5 80 42 ;
        RECT 78.15 42.275 80 42.775 ;
        RECT 78.15 43.05 80 43.55 ;
      LAYER M2 ;
        RECT 78.15 39.95 80 40.45 ;
        RECT 78.15 40.725 80 41.225 ;
        RECT 78.15 41.5 80 42 ;
        RECT 78.15 42.275 80 42.775 ;
        RECT 78.15 43.05 80 43.55 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 77.975 40.25 80 43.25 ;
    END
  END VRES1_B
  PIN VESD3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 24.7745 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 93.505 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 7.05 80 7.55 ;
        RECT 78.15 7.825 80 8.325 ;
        RECT 78.15 8.6 80 9.1 ;
        RECT 78.15 9.375 80 9.875 ;
        RECT 78.15 10.15 80 10.65 ;
      LAYER M2 ;
        RECT 78.15 7.05 80 7.55 ;
        RECT 78.15 7.825 80 8.325 ;
        RECT 78.15 8.6 80 9.1 ;
        RECT 78.15 9.375 80 9.875 ;
        RECT 78.15 10.15 80 10.65 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 77.975 7.35 80 10.35 ;
    END
  END VESD3_B
  PIN VESD2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 21.2495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 96.1675 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.304864 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 21.15 80 21.65 ;
        RECT 78.15 21.925 80 22.425 ;
        RECT 78.15 22.7 80 23.2 ;
        RECT 78.15 23.475 80 23.975 ;
        RECT 78.15 24.25 80 24.75 ;
      LAYER M2 ;
        RECT 78.15 21.15 80 21.65 ;
        RECT 78.15 21.925 80 22.425 ;
        RECT 78.15 22.7 80 23.2 ;
        RECT 78.15 23.475 80 23.975 ;
        RECT 78.15 24.25 80 24.75 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 77.975 21.45 80 24.45 ;
    END
  END VESD2_B
  PIN VRES2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.235 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 22.887 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 85.36 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 7.36 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.304864 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 16.45 80 16.95 ;
        RECT 78.15 17.225 80 17.725 ;
        RECT 78.15 18 80 18.5 ;
        RECT 78.15 18.775 80 19.275 ;
        RECT 78.15 19.55 80 20.05 ;
      LAYER M2 ;
        RECT 78.15 16.45 80 16.95 ;
        RECT 78.15 17.225 80 17.725 ;
        RECT 78.15 18 80 18.5 ;
        RECT 78.15 18.775 80 19.275 ;
        RECT 78.15 19.55 80 20.05 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 77.975 16.75 80 19.75 ;
    END
  END VRES2_B
  PIN VESD1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 42.1975 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 98.0425 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.3392 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 35.25 80 35.75 ;
        RECT 78.15 36.025 80 36.525 ;
        RECT 78.15 36.8 80 37.3 ;
        RECT 78.15 37.575 80 38.075 ;
        RECT 78.15 38.35 80 38.85 ;
      LAYER M2 ;
        RECT 78.15 35.25 80 35.75 ;
        RECT 78.15 36.025 80 36.525 ;
        RECT 78.15 36.8 80 37.3 ;
        RECT 78.15 37.575 80 38.075 ;
        RECT 78.15 38.35 80 38.85 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 77.975 35.55 80 38.55 ;
    END
  END VESD1_B
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_ANACORE_H

MACRO RIIO_EG1D80V_ANAIO_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_ANAIO_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 95.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 567.2075 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 22.385 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 603.245 LAYER IA ;
    ANTENNAPARTIALMETALAREA 294.725 LAYER IB ;
    ANTENNAPARTIALMETALAREA 124.425 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 12.04192 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 7.294848 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 11.54736 LAYER YX ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER XA ;
    ANTENNAPARTIALCUTAREA 4.905824 LAYER A2 ;
    ANTENNADIFFAREA 148.5876 LAYER C4 ;
    ANTENNADIFFAREA 148.5876 LAYER C3 ;
    ANTENNADIFFAREA 148.5876 LAYER C5 ;
    ANTENNADIFFAREA 148.5876 LAYER C6 ;
    ANTENNADIFFAREA 148.5876 LAYER IA ;
    ANTENNADIFFAREA 148.5876 LAYER IB ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN VRES3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 85.987 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 138.78 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.4675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.099 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.747296 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.6144 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.1664 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 44.65 80 45.15 ;
        RECT 78.15 45.425 80 45.925 ;
        RECT 78.15 46.2 80 46.7 ;
        RECT 78.15 46.975 80 47.475 ;
        RECT 78.15 47.75 80 48.25 ;
      LAYER M2 ;
        RECT 78.15 44.65 80 45.15 ;
        RECT 78.15 45.425 80 45.925 ;
        RECT 78.15 46.2 80 46.7 ;
        RECT 78.15 46.975 80 47.475 ;
        RECT 78.15 47.75 80 48.25 ;
      LAYER C1 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 77.975 44.95 80 47.95 ;
    END
  END VRES3_B
  PIN VESD0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 43.4095 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 138.505 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 7.05 80 7.55 ;
        RECT 78.15 7.825 80 8.325 ;
        RECT 78.15 8.6 80 9.1 ;
        RECT 78.15 9.375 80 9.875 ;
        RECT 78.15 10.15 80 10.65 ;
      LAYER M2 ;
        RECT 78.15 7.05 80 7.55 ;
        RECT 78.15 7.825 80 8.325 ;
        RECT 78.15 8.6 80 9.1 ;
        RECT 78.15 9.375 80 9.875 ;
        RECT 78.15 10.15 80 10.65 ;
      LAYER C1 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 77.975 7.35 80 10.35 ;
    END
  END VESD0_B
  PIN VRES0_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.735 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 115.654 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 138.78 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.4675 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.3648 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 11.75 80 12.25 ;
        RECT 78.15 12.525 80 13.025 ;
        RECT 78.15 13.3 80 13.8 ;
        RECT 78.15 14.075 80 14.575 ;
        RECT 78.15 14.85 80 15.35 ;
      LAYER M2 ;
        RECT 78.15 11.75 80 12.25 ;
        RECT 78.15 12.525 80 13.025 ;
        RECT 78.15 13.3 80 13.8 ;
        RECT 78.15 14.075 80 14.575 ;
        RECT 78.15 14.85 80 15.35 ;
      LAYER C1 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 77.975 12.05 80 15.05 ;
    END
  END VRES0_B
  PIN VRES1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.235 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 41.522 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 132.235 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 7.36 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.204192 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 16.45 80 16.95 ;
        RECT 78.15 17.225 80 17.725 ;
        RECT 78.15 18 80 18.5 ;
        RECT 78.15 18.775 80 19.275 ;
        RECT 78.15 19.55 80 20.05 ;
      LAYER M2 ;
        RECT 78.15 16.45 80 16.95 ;
        RECT 78.15 17.225 80 17.725 ;
        RECT 78.15 18 80 18.5 ;
        RECT 78.15 18.775 80 19.275 ;
        RECT 78.15 19.55 80 20.05 ;
      LAYER C1 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 77.975 16.75 80 19.75 ;
    END
  END VRES1_B
  PIN VESD3_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 43.4095 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 138.505 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 63.1925 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 49.35 80 49.85 ;
        RECT 78.15 50.125 80 50.625 ;
        RECT 78.15 50.9 80 51.4 ;
        RECT 78.15 51.675 80 52.175 ;
        RECT 78.15 52.45 80 52.95 ;
      LAYER M2 ;
        RECT 78.15 49.35 80 49.85 ;
        RECT 78.15 50.125 80 50.625 ;
        RECT 78.15 50.9 80 51.4 ;
        RECT 78.15 51.675 80 52.175 ;
        RECT 78.15 52.45 80 52.95 ;
      LAYER C1 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 77.975 49.65 80 52.65 ;
    END
  END VESD3_B
  PIN VESD2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 60.1975 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 143.805 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.3392 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 35.25 80 35.75 ;
        RECT 78.15 36.025 80 36.525 ;
        RECT 78.15 36.8 80 37.3 ;
        RECT 78.15 37.575 80 38.075 ;
        RECT 78.15 38.35 80 38.85 ;
      LAYER M2 ;
        RECT 78.15 35.25 80 35.75 ;
        RECT 78.15 36.025 80 36.525 ;
        RECT 78.15 36.8 80 37.3 ;
        RECT 78.15 37.575 80 38.075 ;
        RECT 78.15 38.35 80 38.85 ;
      LAYER C1 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 77.975 35.55 80 38.55 ;
    END
  END VESD2_B
  PIN VRES2_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.235 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 41.522 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 132.235 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 39.95 80 40.45 ;
        RECT 78.15 40.725 80 41.225 ;
        RECT 78.15 41.5 80 42 ;
        RECT 78.15 42.275 80 42.775 ;
        RECT 78.15 43.05 80 43.55 ;
      LAYER M2 ;
        RECT 78.15 39.95 80 40.45 ;
        RECT 78.15 40.725 80 41.225 ;
        RECT 78.15 41.5 80 42 ;
        RECT 78.15 42.275 80 42.775 ;
        RECT 78.15 43.05 80 43.55 ;
      LAYER C1 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 77.975 40.25 80 43.25 ;
    END
  END VRES2_B
  PIN VESD1_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 39.8845 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 143.805 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 32.36 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 13.61 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 56.9225 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER IA ;
    ANTENNAPARTIALMETALAREA 1.11 LAYER IB ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 1.444256 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 0.1856 LAYER AY ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 1.80048 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 0.607904 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER YX ;
    ANTENNAPARTIALCUTAREA 1.04976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 0.416 LAYER V1 ;
    ANTENNADIFFAREA 20.425 LAYER C3 ;
    ANTENNADIFFAREA 20.425 LAYER C2 ;
    ANTENNADIFFAREA 20.425 LAYER C4 ;
    ANTENNADIFFAREA 20.425 LAYER C5 ;
    ANTENNADIFFAREA 20.425 LAYER C6 ;
    ANTENNADIFFAREA 20.425 LAYER IA ;
    ANTENNADIFFAREA 20.425 LAYER IB ;
    ANTENNADIFFAREA 20.425 LAYER C1 ;
    PORT
      LAYER M1 ;
        RECT 78.15 21.15 80 21.65 ;
        RECT 78.15 21.925 80 22.425 ;
        RECT 78.15 22.7 80 23.2 ;
        RECT 78.15 23.475 80 23.975 ;
        RECT 78.15 24.25 80 24.75 ;
      LAYER M2 ;
        RECT 78.15 21.15 80 21.65 ;
        RECT 78.15 21.925 80 22.425 ;
        RECT 78.15 22.7 80 23.2 ;
        RECT 78.15 23.475 80 23.975 ;
        RECT 78.15 24.25 80 24.75 ;
      LAYER C1 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 77.975 21.45 80 24.45 ;
    END
  END VESD1_B
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_ANAIO_H

MACRO RIIO_EG1D80V_BIASPAD_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_BIASPAD_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.25 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 46.875 LAYER C5 ;
    ANTENNAPARTIALCUTAREA 0.894432 LAYER A4 ;
    ANTENNADIFFAREA 3.608 LAYER C4 ;
    ANTENNADIFFAREA 3.608 LAYER C5 ;
    NETEXPR "vbias VBIAS!" ;
    PORT
      LAYER C4 ;
        RECT 39.575 0 40.825 60 ;
    END
  END VBIAS
  PIN PAD_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 370.645 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 198.8 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 381.9382 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 529.985 LAYER IA ;
    ANTENNAPARTIALMETALAREA 294.725 LAYER IB ;
    ANTENNAPARTIALMETALAREA 244.78 LAYER C2 ;
    ANTENNAPARTIALCUTAREA 11.434016 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 13.257728 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 4.905824 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 31.4928 LAYER YX ;
    ANTENNAPARTIALCUTAREA 27.713664 LAYER XA ;
    ANTENNAPARTIALCUTAREA 6.055808 LAYER A2 ;
    ANTENNADIFFAREA 148.5876 LAYER C4 ;
    ANTENNADIFFAREA 148.5876 LAYER C3 ;
    ANTENNADIFFAREA 148.5876 LAYER C5 ;
    ANTENNADIFFAREA 148.5876 LAYER C6 ;
    ANTENNADIFFAREA 148.5876 LAYER IA ;
    ANTENNADIFFAREA 148.5876 LAYER IB ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT -0.001 2.35 1.849 5.95 ;
        RECT -0.001 7.05 1.849 10.65 ;
        RECT -0.001 11.75 1.849 15.35 ;
        RECT -0.001 16.45 1.849 20.05 ;
        RECT -0.001 21.15 1.849 24.75 ;
        RECT -0.001 25.85 1.849 29.45 ;
        RECT -0.001 30.55 1.849 34.15 ;
        RECT -0.001 35.25 1.849 38.85 ;
        RECT -0.001 39.95 1.849 43.55 ;
        RECT -0.001 44.65 1.849 48.25 ;
        RECT -0.001 49.35 1.849 52.95 ;
        RECT -0.001 54.05 1.849 57.65 ;
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
  END PAD_B
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_BIASPAD_H

MACRO RIIO_EG1D80V_CUTB2B_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTB2B_H 0 0 ;
  SIZE 80 BY 16 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_l VSS_L!" ;
    PORT
      LAYER IB ;
        RECT 59.35 10 62.95 16 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 10 77.05 16 ;
    END
  END VSS_L
  PIN VSS_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_r VSS_R!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 6 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 6 ;
    END
  END VSS_R
  PIN VSSIO_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_l VSSIO_L!" ;
    PORT
      LAYER IB ;
        RECT 3.67 10 6.55 16 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 10 20.65 16 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 10 30.05 16 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 10 44.15 16 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 10 48.85 16 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 10 58.25 16 ;
    END
  END VSSIO_L
  PIN VSSIO_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_r VSSIO_R!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 6 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 6 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 6 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 6 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 6 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 6 ;
    END
  END VSSIO_R
  OBS
    LAYER CA ;
      RECT 0 0 80 16 ;
    LAYER M1 ;
      RECT 0 0 80 16 ;
    LAYER V1 ;
      RECT 0 0 80 16 ;
    LAYER M2 ;
      RECT 0 0 80 16 ;
    LAYER A1 ;
      RECT 0 0 80 16 ;
    LAYER C2 ;
      RECT 0 0 80 16 ;
    LAYER IA ;
      RECT 0 0 80 16 ;
    LAYER XA ;
      RECT 0 0 80 16 ;
    LAYER YX ;
      RECT 0 0 80 16 ;
    LAYER IB ;
      RECT 0 0 80 16 ;
    LAYER CB ;
      RECT 0 0 80 16 ;
    LAYER AY ;
      RECT 0 0 80 16 ;
    LAYER C1 ;
      RECT 0 0 80 16 ;
    LAYER C5 ;
      RECT 0 0 80 16 ;
    LAYER C4 ;
      RECT 0 0 80 16 ;
    LAYER C3 ;
      RECT 0 0 80 16 ;
    LAYER A5 ;
      RECT 0 0 80 16 ;
    LAYER A4 ;
      RECT 0 0 80 16 ;
    LAYER A3 ;
      RECT 0 0 80 16 ;
    LAYER A2 ;
      RECT 0 0 80 16 ;
    LAYER C6 ;
      RECT 0 0 80 16 ;
  END
END RIIO_EG1D80V_CUTB2B_H

MACRO RIIO_EG1D80V_CUTBIAS_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTBIAS_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 4 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 4 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 4 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 4 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 4 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 4 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 4 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 4 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTBIAS_H

MACRO RIIO_EG1D80V_CUTCOREB2B_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCOREB2B_H 0 0 ;
  SIZE 80 BY 16 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 16 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 16 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 16 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 16 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 16 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 16 ;
    END
  END VSSIO
  PIN VSS_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_l VSS_L!" ;
    PORT
      LAYER IB ;
        RECT 59.35 10 62.95 16 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 10 77.05 16 ;
    END
  END VSS_L
  PIN VSS_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_r VSS_R!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 6 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 6 ;
    END
  END VSS_R
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 16 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 16 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 16 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 16 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 16 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 16 ;
    LAYER M1 ;
      RECT 0 0 80 16 ;
    LAYER V1 ;
      RECT 0 0 80 16 ;
    LAYER M2 ;
      RECT 0 0 80 16 ;
    LAYER A1 ;
      RECT 0 0 80 16 ;
    LAYER C2 ;
      RECT 0 0 80 16 ;
    LAYER IA ;
      RECT 0 0 80 16 ;
    LAYER XA ;
      RECT 0 0 80 16 ;
    LAYER YX ;
      RECT 0 0 80 16 ;
    LAYER IB ;
      RECT 0 0 80 16 ;
    LAYER CB ;
      RECT 0 0 80 16 ;
    LAYER AY ;
      RECT 0 0 80 16 ;
    LAYER C1 ;
      RECT 0 0 80 16 ;
    LAYER C5 ;
      RECT 0 0 80 16 ;
    LAYER C4 ;
      RECT 0 0 80 16 ;
    LAYER C3 ;
      RECT 0 0 80 16 ;
    LAYER A5 ;
      RECT 0 0 80 16 ;
    LAYER A4 ;
      RECT 0 0 80 16 ;
    LAYER A3 ;
      RECT 0 0 80 16 ;
    LAYER A2 ;
      RECT 0 0 80 16 ;
    LAYER C6 ;
      RECT 0 0 80 16 ;
  END
END RIIO_EG1D80V_CUTCOREB2B_H

MACRO RIIO_EG1D80V_CUTCOREPWR_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCOREPWR_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 4 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 4 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 4 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 4 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 4 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 4 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 4 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 4 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTCOREPWR_H

MACRO RIIO_EG1D80V_CUTCORE_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTCORE_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 4 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 4 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 4 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 4 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 4 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 4 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 4 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTCORE_H

MACRO RIIO_EG1D80V_CUTIOB2B_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIOB2B_H 0 0 ;
  SIZE 80 BY 16 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 16 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 16 ;
    END
  END VSS
  PIN VSSIO_L
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_l VSSIO_L!" ;
    PORT
      LAYER IB ;
        RECT 3.67 10 6.55 16 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 10 20.65 16 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 10 30.05 16 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 10 44.15 16 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 10 48.85 16 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 10 58.25 16 ;
    END
  END VSSIO_L
  PIN VSSIO_R
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_r VSSIO_R!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 6 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 6 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 6 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 6 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 6 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 6 ;
    END
  END VSSIO_R
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 16 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 16 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 16 ;
    LAYER M1 ;
      RECT 0 0 80 16 ;
    LAYER V1 ;
      RECT 0 0 80 16 ;
    LAYER M2 ;
      RECT 0 0 80 16 ;
    LAYER A1 ;
      RECT 0 0 80 16 ;
    LAYER C2 ;
      RECT 0 0 80 16 ;
    LAYER IA ;
      RECT 0 0 80 16 ;
    LAYER XA ;
      RECT 0 0 80 16 ;
    LAYER YX ;
      RECT 0 0 80 16 ;
    LAYER IB ;
      RECT 0 0 80 16 ;
    LAYER CB ;
      RECT 0 0 80 16 ;
    LAYER AY ;
      RECT 0 0 80 16 ;
    LAYER C1 ;
      RECT 0 0 80 16 ;
    LAYER C5 ;
      RECT 0 0 80 16 ;
    LAYER C4 ;
      RECT 0 0 80 16 ;
    LAYER C3 ;
      RECT 0 0 80 16 ;
    LAYER A5 ;
      RECT 0 0 80 16 ;
    LAYER A4 ;
      RECT 0 0 80 16 ;
    LAYER A3 ;
      RECT 0 0 80 16 ;
    LAYER A2 ;
      RECT 0 0 80 16 ;
    LAYER C6 ;
      RECT 0 0 80 16 ;
  END
END RIIO_EG1D80V_CUTIOB2B_H

MACRO RIIO_EG1D80V_CUTIOPWR_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIOPWR_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 4 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 4 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 4 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 4 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 4 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTIOPWR_H

MACRO RIIO_EG1D80V_CUTIO_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTIO_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 4 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTIO_H

MACRO RIIO_EG1D80V_CUTPWR_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUTPWR_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 4 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 4 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 4 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 4 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 4 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUTPWR_H

MACRO RIIO_EG1D80V_CUT_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_CUT_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_CUT_H

MACRO RIIO_EG1D80V_FILL16B2B_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL16B2B_H 0 0 ;
  SIZE 80 BY 16 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 16 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 16 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 16 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 16 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 16 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 16 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 16 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 16 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 16 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 16 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 16 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 16 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 16 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 16 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 16 ;
    LAYER M1 ;
      RECT 0 0 80 16 ;
    LAYER V1 ;
      RECT 0 0 80 16 ;
    LAYER M2 ;
      RECT 0 0 80 16 ;
    LAYER A1 ;
      RECT 0 0 80 16 ;
    LAYER C2 ;
      RECT 0 0 80 16 ;
    LAYER IA ;
      RECT 0 0 80 16 ;
    LAYER XA ;
      RECT 0 0 80 16 ;
    LAYER YX ;
      RECT 0 0 80 16 ;
    LAYER IB ;
      RECT 0 0 80 16 ;
    LAYER CB ;
      RECT 0 0 80 16 ;
    LAYER AY ;
      RECT 0 0 80 16 ;
    LAYER C1 ;
      RECT 0 0 80 16 ;
    LAYER C5 ;
      RECT 0 0 80 16 ;
    LAYER C4 ;
      RECT 0 0 80 16 ;
    LAYER C3 ;
      RECT 0 0 80 16 ;
    LAYER A5 ;
      RECT 0 0 80 16 ;
    LAYER A4 ;
      RECT 0 0 80 16 ;
    LAYER A3 ;
      RECT 0 0 80 16 ;
    LAYER A2 ;
      RECT 0 0 80 16 ;
    LAYER C6 ;
      RECT 0 0 80 16 ;
  END
END RIIO_EG1D80V_FILL16B2B_H

MACRO RIIO_EG1D80V_FILL16_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL16_H 0 0 ;
  SIZE 80 BY 16 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 16 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 16 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 16 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 16 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 16 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 16 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 16 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 16 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 16 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 16 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 16 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 16 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 16 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 16 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 16 ;
    LAYER M1 ;
      RECT 0 0 80 16 ;
    LAYER V1 ;
      RECT 0 0 80 16 ;
    LAYER M2 ;
      RECT 0 0 80 16 ;
    LAYER A1 ;
      RECT 0 0 80 16 ;
    LAYER C2 ;
      RECT 0 0 80 16 ;
    LAYER IA ;
      RECT 0 0 80 16 ;
    LAYER XA ;
      RECT 0 0 80 16 ;
    LAYER YX ;
      RECT 0 0 80 16 ;
    LAYER IB ;
      RECT 0 0 80 16 ;
    LAYER CB ;
      RECT 0 0 80 16 ;
    LAYER AY ;
      RECT 0 0 80 16 ;
    LAYER C1 ;
      RECT 0 0 80 16 ;
    LAYER C5 ;
      RECT 0 0 80 16 ;
    LAYER C4 ;
      RECT 0 0 80 16 ;
    LAYER C3 ;
      RECT 0 0 80 16 ;
    LAYER A5 ;
      RECT 0 0 80 16 ;
    LAYER A4 ;
      RECT 0 0 80 16 ;
    LAYER A3 ;
      RECT 0 0 80 16 ;
    LAYER A2 ;
      RECT 0 0 80 16 ;
    LAYER C6 ;
      RECT 0 0 80 16 ;
  END
END RIIO_EG1D80V_FILL16_H

MACRO RIIO_EG1D80V_FILL1_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL1_H 0 0 ;
  SIZE 80 BY 1 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 1 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 1 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 1 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 1 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 1 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 1 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 1 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 1 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 1 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 1 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 1 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 1 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 1 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 1 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 1 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 1 ;
    LAYER M1 ;
      RECT 0 0 80 1 ;
    LAYER V1 ;
      RECT 0 0 80 1 ;
    LAYER M2 ;
      RECT 0 0 80 1 ;
    LAYER A1 ;
      RECT 0 0 80 1 ;
    LAYER C2 ;
      RECT 0 0 80 1 ;
    LAYER IA ;
      RECT 0 0 80 1 ;
    LAYER XA ;
      RECT 0 0 80 1 ;
    LAYER YX ;
      RECT 0 0 80 1 ;
    LAYER IB ;
      RECT 0 0 80 1 ;
    LAYER CB ;
      RECT 0 0 80 1 ;
    LAYER AY ;
      RECT 0 0 80 1 ;
    LAYER C1 ;
      RECT 0 0 80 1 ;
    LAYER C5 ;
      RECT 0 0 80 1 ;
    LAYER C4 ;
      RECT 0 0 80 1 ;
    LAYER C3 ;
      RECT 0 0 80 1 ;
    LAYER A5 ;
      RECT 0 0 80 1 ;
    LAYER A4 ;
      RECT 0 0 80 1 ;
    LAYER A3 ;
      RECT 0 0 80 1 ;
    LAYER A2 ;
      RECT 0 0 80 1 ;
    LAYER C6 ;
      RECT 0 0 80 1 ;
  END
END RIIO_EG1D80V_FILL1_H

MACRO RIIO_EG1D80V_FILL2_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL2_H 0 0 ;
  SIZE 80 BY 2 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 2 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 2 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 2 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 2 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 2 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 2 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 2 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 2 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 2 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 2 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 2 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 2 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 2 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 2 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 2 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 80 2 ;
    LAYER M1 ;
      RECT 0 0 80 2 ;
    LAYER V1 ;
      RECT 0 0 80 2 ;
    LAYER M2 ;
      RECT 0 0 80 2 ;
    LAYER A1 ;
      RECT 0 0 80 2 ;
    LAYER C2 ;
      RECT 0 0 80 2 ;
    LAYER IA ;
      RECT 0 0 80 2 ;
    LAYER XA ;
      RECT 0 0 80 2 ;
    LAYER YX ;
      RECT 0 0 80 2 ;
    LAYER IB ;
      RECT 0 0 80 2 ;
    LAYER CB ;
      RECT 0 0 80 2 ;
    LAYER AY ;
      RECT 0 0 80 2 ;
    LAYER C1 ;
      RECT 0 0 80 2 ;
    LAYER C5 ;
      RECT 0 0 80 2 ;
    LAYER C4 ;
      RECT 0 0 80 2 ;
    LAYER C3 ;
      RECT 0 0 80 2 ;
    LAYER A5 ;
      RECT 0 0 80 2 ;
    LAYER A4 ;
      RECT 0 0 80 2 ;
    LAYER A3 ;
      RECT 0 0 80 2 ;
    LAYER A2 ;
      RECT 0 0 80 2 ;
    LAYER C6 ;
      RECT 0 0 80 2 ;
  END
END RIIO_EG1D80V_FILL2_H

MACRO RIIO_EG1D80V_FILL32_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL32_H 0 0 ;
  SIZE 80 BY 32 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 32 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 32 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 32 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 32 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 32 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 32 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 32 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 32 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 32 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 32 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 32 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 32 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 32 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 32 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 32 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 80 32 ;
    LAYER M1 ;
      RECT 0 0 80 32 ;
    LAYER V1 ;
      RECT 0 0 80 32 ;
    LAYER M2 ;
      RECT 0 0 80 32 ;
    LAYER A1 ;
      RECT 0 0 80 32 ;
    LAYER C2 ;
      RECT 0 0 80 32 ;
    LAYER IA ;
      RECT 0 0 80 32 ;
    LAYER XA ;
      RECT 0 0 80 32 ;
    LAYER YX ;
      RECT 0 0 80 32 ;
    LAYER IB ;
      RECT 0 0 80 32 ;
    LAYER CB ;
      RECT 0 0 80 32 ;
    LAYER AY ;
      RECT 0 0 80 32 ;
    LAYER C1 ;
      RECT 0 0 80 32 ;
    LAYER C5 ;
      RECT 0 0 80 32 ;
    LAYER C4 ;
      RECT 0 0 80 32 ;
    LAYER C3 ;
      RECT 0 0 80 32 ;
    LAYER A5 ;
      RECT 0 0 80 32 ;
    LAYER A4 ;
      RECT 0 0 80 32 ;
    LAYER A3 ;
      RECT 0 0 80 32 ;
    LAYER A2 ;
      RECT 0 0 80 32 ;
    LAYER C6 ;
      RECT 0 0 80 32 ;
  END
END RIIO_EG1D80V_FILL32_H

MACRO RIIO_EG1D80V_FILL4_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL4_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 4 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 4 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 4 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 4 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 4 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 4 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 4 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 4 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_FILL4_H

MACRO RIIO_EG1D80V_FILL8_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_FILL8_H 0 0 ;
  SIZE 80 BY 8 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 8 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 8 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 8 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 8 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 8 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 8 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 8 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 8 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 8 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 8 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 8 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 8 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 8 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 8 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 8 ;
    LAYER M1 ;
      RECT 0 0 80 8 ;
    LAYER V1 ;
      RECT 0 0 80 8 ;
    LAYER M2 ;
      RECT 0 0 80 8 ;
    LAYER A1 ;
      RECT 0 0 80 8 ;
    LAYER C2 ;
      RECT 0 0 80 8 ;
    LAYER IA ;
      RECT 0 0 80 8 ;
    LAYER XA ;
      RECT 0 0 80 8 ;
    LAYER YX ;
      RECT 0 0 80 8 ;
    LAYER IB ;
      RECT 0 0 80 8 ;
    LAYER CB ;
      RECT 0 0 80 8 ;
    LAYER AY ;
      RECT 0 0 80 8 ;
    LAYER C1 ;
      RECT 0 0 80 8 ;
    LAYER C5 ;
      RECT 0 0 80 8 ;
    LAYER C4 ;
      RECT 0 0 80 8 ;
    LAYER C3 ;
      RECT 0 0 80 8 ;
    LAYER A5 ;
      RECT 0 0 80 8 ;
    LAYER A4 ;
      RECT 0 0 80 8 ;
    LAYER A3 ;
      RECT 0 0 80 8 ;
    LAYER A2 ;
      RECT 0 0 80 8 ;
    LAYER C6 ;
      RECT 0 0 80 8 ;
  END
END RIIO_EG1D80V_FILL8_H

MACRO RIIO_EG1D80V_POR_IO_V1D0_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_POR_IO_V1D0_H 0 0 ;
  SIZE 80 BY 8 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER C3 ;
        RECT 37.075 0 39.575 8 ;
    END
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 8 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 8 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 8 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 8 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 8 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 8 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 8 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 8 ;
      LAYER C3 ;
        RECT 70.825 0 73.325 8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 8 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 8 ;
      LAYER C3 ;
        RECT 74.575 0 77.075 8 ;
    END
  END VSS
  PIN VDDIO_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio_por VDDIO_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 33.325 2.625 80 3.125 ;
    END
  END VDDIO_POR
  PIN POR_N_CORE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3375 LAYER C2 ;
    ANTENNADIFFAREA 0.2453 LAYER C2 ;
    PORT
      LAYER C2 ;
        RECT 79.5 5.625 80 6.125 ;
    END
  END POR_N_CORE_O
  PIN VDD_POR
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd_por VDD_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 70.825 4.125 80 4.625 ;
    END
  END VDD_POR
  PIN VSSIO_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio_por VSSIO_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 33.325 1.875 80 2.375 ;
    END
  END VSSIO_POR
  PIN VSS_POR
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss_por VSS_POR!" ;
    PORT
      CLASS CORE ;
      LAYER C2 ;
        RECT 70.825 4.875 80 5.375 ;
    END
  END VSS_POR
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 8 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 8 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 8 ;
      LAYER C3 ;
        RECT 33.325 0 35.825 8 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 8 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 8 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 8 ;
    LAYER M1 ;
      RECT 0 0 80 8 ;
    LAYER V1 ;
      RECT 0 0 80 8 ;
    LAYER M2 ;
      RECT 0 0 80 8 ;
    LAYER A1 ;
      RECT 0 0 80 8 ;
    LAYER C2 ;
      RECT 0 0 80 8 ;
    LAYER IA ;
      RECT 0 0 80 8 ;
    LAYER XA ;
      RECT 0 0 80 8 ;
    LAYER YX ;
      RECT 0 0 80 8 ;
    LAYER IB ;
      RECT 0 0 80 8 ;
    LAYER CB ;
      RECT 0 0 80 8 ;
    LAYER AY ;
      RECT 0 0 80 8 ;
    LAYER C1 ;
      RECT 0 0 80 8 ;
    LAYER C5 ;
      RECT 0 0 80 8 ;
    LAYER C4 ;
      RECT 0 0 80 8 ;
    LAYER C3 ;
      RECT 0 0 80 8 ;
    LAYER A5 ;
      RECT 0 0 80 8 ;
    LAYER A4 ;
      RECT 0 0 80 8 ;
    LAYER A3 ;
      RECT 0 0 80 8 ;
    LAYER A2 ;
      RECT 0 0 80 8 ;
    LAYER C6 ;
      RECT 0 0 80 8 ;
  END
END RIIO_EG1D80V_POR_IO_V1D0_H

MACRO RIIO_EG1D80V_RAILSHORT_GND_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_GND_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 4 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 4 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 4 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 4 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 4 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 4 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 4 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 4 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 4 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_RAILSHORT_GND_H

MACRO RIIO_EG1D80V_RAILSHORT_PG_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_PG_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 4 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 4 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 4 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 4 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 4 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 4 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 4 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 4 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_RAILSHORT_PG_H

MACRO RIIO_EG1D80V_RAILSHORT_PWR_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_RAILSHORT_PWR_H 0 0 ;
  SIZE 80 BY 4 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 4 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 4 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 4 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 4 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 4 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 4 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 4 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 4 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 4 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 4 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 4 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 4 ;
    LAYER M1 ;
      RECT 0 0 80 4 ;
    LAYER V1 ;
      RECT 0 0 80 4 ;
    LAYER M2 ;
      RECT 0 0 80 4 ;
    LAYER A1 ;
      RECT 0 0 80 4 ;
    LAYER C2 ;
      RECT 0 0 80 4 ;
    LAYER IA ;
      RECT 0 0 80 4 ;
    LAYER XA ;
      RECT 0 0 80 4 ;
    LAYER YX ;
      RECT 0 0 80 4 ;
    LAYER IB ;
      RECT 0 0 80 4 ;
    LAYER CB ;
      RECT 0 0 80 4 ;
    LAYER AY ;
      RECT 0 0 80 4 ;
    LAYER C1 ;
      RECT 0 0 80 4 ;
    LAYER C5 ;
      RECT 0 0 80 4 ;
    LAYER C4 ;
      RECT 0 0 80 4 ;
    LAYER C3 ;
      RECT 0 0 80 4 ;
    LAYER A5 ;
      RECT 0 0 80 4 ;
    LAYER A4 ;
      RECT 0 0 80 4 ;
    LAYER A3 ;
      RECT 0 0 80 4 ;
    LAYER A2 ;
      RECT 0 0 80 4 ;
    LAYER C6 ;
      RECT 0 0 80 4 ;
  END
END RIIO_EG1D80V_RAILSHORT_PWR_H

MACRO RIIO_EG1D80V_VDD04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDD04_H

MACRO RIIO_EG1D80V_VDDIOX_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDIOX_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIOX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddiox VDDIOX!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDDIOX
  PIN VSSIOX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssiox VSSIOX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C1 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER M2 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
  END VSSIOX
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDIOX_H

MACRO RIIO_EG1D80V_VDDIO_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDIO_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDIO_H

MACRO RIIO_EG1D80V_VDDQ04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSQ
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDDQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDQ04_H

MACRO RIIO_EG1D80V_VDDQ_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSQ
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDDQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDQ_HVT_H

MACRO RIIO_EG1D80V_VDDQ_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDQ_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSQ
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDDQ
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDQ_RVT_H

MACRO RIIO_EG1D80V_VDDX04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 47.5 80 50 ;
      LAYER M2 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER C1 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 17.5 80 20 ;
      LAYER M2 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER C1 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
  END VSSX
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDX04_H

MACRO RIIO_EG1D80V_VDDX_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C1 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER M2 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDX_HVT_H

MACRO RIIO_EG1D80V_VDDX_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDDX_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C1 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER M2 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDDX_RVT_H

MACRO RIIO_EG1D80V_VDD_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 54.393 79.958 57.393 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 49.693 79.958 52.693 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 44.993 79.958 47.993 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 40.293 79.958 43.293 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 35.593 79.958 38.593 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 30.893 79.958 33.893 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 26.193 79.958 29.193 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 21.493 79.958 24.493 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 16.793 79.958 19.793 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 12.093 79.958 15.093 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 7.393 79.958 10.393 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 2.693 79.958 5.693 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT -0.042 54.093 1.808 57.693 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT -0.042 49.393 1.808 52.993 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT -0.042 44.693 1.808 48.293 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT -0.042 39.993 1.808 43.593 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT -0.042 35.293 1.808 38.893 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT -0.042 30.593 1.808 34.193 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT -0.042 25.893 1.808 29.493 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT -0.042 21.193 1.808 24.793 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT -0.042 16.493 1.808 20.093 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT -0.042 11.793 1.808 15.393 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT -0.042 7.093 1.808 10.693 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT -0.042 2.393 1.808 5.993 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDD_HVT_H

MACRO RIIO_EG1D80V_VDD_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VDD_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 54.393 79.958 57.393 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 49.693 79.958 52.693 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 44.993 79.958 47.993 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 40.293 79.958 43.293 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 35.593 79.958 38.593 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 30.893 79.958 33.893 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 26.193 79.958 29.193 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 21.493 79.958 24.493 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 16.793 79.958 19.793 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 12.093 79.958 15.093 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 7.393 79.958 10.393 ;
    END
    PORT
      LAYER C6 ;
        RECT 78.108 2.693 79.958 5.693 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT -0.042 54.093 1.808 57.693 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT -0.042 49.393 1.808 52.993 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT -0.042 44.693 1.808 48.293 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT -0.042 39.993 1.808 43.593 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT -0.042 35.293 1.808 38.893 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT -0.042 30.593 1.808 34.193 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT -0.042 25.893 1.808 29.493 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT -0.042 21.193 1.808 24.793 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT -0.042 16.493 1.808 20.093 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT -0.042 11.793 1.808 15.393 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT -0.042 7.093 1.808 10.693 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT -0.042 2.393 1.808 5.993 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VDD_RVT_H

MACRO RIIO_EG1D80V_VNWINT_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNWINT_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.103 1.85 57.703 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.403 1.85 53.003 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.703 1.85 48.303 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 40.003 1.85 43.603 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.303 1.85 38.903 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.603 1.85 34.203 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.903 1.85 29.503 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.203 1.85 24.803 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.503 1.85 20.103 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.803 1.85 15.403 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.103 1.85 10.703 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.403 1.85 6.003 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.403 80 57.403 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.703 80 52.703 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 45.003 80 48.003 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.303 80 43.303 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.603 80 38.603 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.903 80 33.903 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.203 80 29.203 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.503 80 24.503 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.803 80 19.803 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.103 80 15.103 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.403 80 10.403 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.703 80 5.703 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VNWINT_HVT_H

MACRO RIIO_EG1D80V_VNWINT_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNWINT_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.103 1.85 57.703 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.403 1.85 53.003 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.703 1.85 48.303 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 40.003 1.85 43.603 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.303 1.85 38.903 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.603 1.85 34.203 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.903 1.85 29.503 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.203 1.85 24.803 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.503 1.85 20.103 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.803 1.85 15.403 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.103 1.85 10.703 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.403 1.85 6.003 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.403 80 57.403 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.703 80 52.703 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 45.003 80 48.003 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.303 80 43.303 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.603 80 38.603 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.903 80 33.903 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.203 80 29.203 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.503 80 24.503 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.803 80 19.803 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.103 80 15.103 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.403 80 10.403 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.703 80 5.703 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VNWINT_RVT_H

MACRO RIIO_EG1D80V_VNW_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VNW_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vnw VNW!" ;
    PORT
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.103 1.85 57.703 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.403 1.85 53.003 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.703 1.85 48.303 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 40.003 1.85 43.603 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.303 1.85 38.903 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.603 1.85 34.203 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.903 1.85 29.503 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.203 1.85 24.803 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.503 1.85 20.103 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.803 1.85 15.403 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.103 1.85 10.703 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.403 1.85 6.003 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.403 80 57.403 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.703 80 52.703 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 45.003 80 48.003 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.303 80 43.303 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.603 80 38.603 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.903 80 33.903 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.203 80 29.203 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.503 80 24.503 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.803 80 19.803 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.103 80 15.103 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.403 80 10.403 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.703 80 5.703 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VNW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VNW_H

MACRO RIIO_EG1D80V_VPWINT_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPWINT_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VPWINT_HVT_H

MACRO RIIO_EG1D80V_VPWINT_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPWINT_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VPWINT_RVT_H

MACRO RIIO_EG1D80V_VPW_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VPW_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vpw VPW!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VPW
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VPW_H

MACRO RIIO_EG1D80V_VSS04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSS04_H

MACRO RIIO_EG1D80V_VSSIOX_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSIOX_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VSSIOX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssiox VSSIOX!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C1 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER M2 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSSIOX
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIOX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddiox VDDIOX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.153 44.95 80.003 47.95 ;
      LAYER C6 ;
        RECT 78.153 44.95 80.003 47.95 ;
      LAYER C5 ;
        RECT 78.153 44.95 80.003 47.95 ;
      LAYER C4 ;
        RECT 78.153 44.95 80.003 47.95 ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER IB ;
        RECT 78.153 44.95 80.003 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.153 40.25 80.003 43.25 ;
      LAYER C6 ;
        RECT 78.153 40.25 80.003 43.25 ;
      LAYER C5 ;
        RECT 78.153 40.25 80.003 43.25 ;
      LAYER C4 ;
        RECT 78.153 40.25 80.003 43.25 ;
      LAYER IB ;
        RECT 78.153 40.25 80.003 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.153 16.75 80.003 19.75 ;
      LAYER C6 ;
        RECT 78.153 16.75 80.003 19.75 ;
      LAYER C5 ;
        RECT 78.153 16.75 80.003 19.75 ;
      LAYER C4 ;
        RECT 78.153 16.75 80.003 19.75 ;
      LAYER IB ;
        RECT 78.153 16.75 80.003 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.153 12.05 80.003 15.05 ;
      LAYER C6 ;
        RECT 78.153 12.05 80.003 15.05 ;
      LAYER C5 ;
        RECT 78.153 12.05 80.003 15.05 ;
      LAYER C4 ;
        RECT 78.153 12.05 80.003 15.05 ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER IB ;
        RECT 78.153 12.05 80.003 15.05 ;
    END
  END VDDIOX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSIOX_H

MACRO RIIO_EG1D80V_VSSIO_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSIO_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSSIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSIO_H

MACRO RIIO_EG1D80V_VSSQ04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDQ
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSQ04_H

MACRO RIIO_EG1D80V_VSSQ_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDQ
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSQ_HVT_H

MACRO RIIO_EG1D80V_VSSQ_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSQ_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VDDQ
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddq VDDQ!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDQ
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VSSQ
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssq VSSQ!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSSQ
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSQ_RVT_H

MACRO RIIO_EG1D80V_VSSX04_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX04_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 17.5 80 20 ;
      LAYER M2 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER C1 ;
        RECT 79.19 17.338 80 20.163 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 47.5 80 50 ;
      LAYER M2 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER C1 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSSX
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSX04_H

MACRO RIIO_EG1D80V_VSSX_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C1 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER M2 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSX_HVT_H

MACRO RIIO_EG1D80V_VSSX_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSSX_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSSX
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssx VSSX!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C2 ;
        RECT 78.15 40 80 42.5 ;
      LAYER C1 ;
        RECT 79.19 39.838 80 42.663 ;
      LAYER M2 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
      LAYER M1 ;
        RECT 79.19 39.838 80 40.338 ;
        RECT 79.19 40.613 80 41.113 ;
        RECT 79.19 41.388 80 41.888 ;
        RECT 79.19 42.163 80 42.663 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C2 ;
        RECT 78.15 17.5 80 20 ;
      LAYER C1 ;
        RECT 79.19 17.338 80 20.163 ;
      LAYER M2 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
      LAYER M1 ;
        RECT 79.19 17.338 80 17.838 ;
        RECT 79.19 18.113 80 18.613 ;
        RECT 79.19 18.888 80 19.388 ;
        RECT 79.19 19.663 80 20.163 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C2 ;
        RECT 78.15 47.5 80 50 ;
      LAYER C1 ;
        RECT 79.19 47.338 80 50.163 ;
      LAYER M2 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER M1 ;
        RECT 79.19 47.338 80 47.838 ;
        RECT 79.19 48.113 80 48.613 ;
        RECT 79.19 48.888 80 49.388 ;
        RECT 79.19 49.663 80 50.163 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C2 ;
        RECT 78.15 32.5 80 35 ;
      LAYER C1 ;
        RECT 79.19 32.338 80 35.163 ;
      LAYER M2 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER M1 ;
        RECT 79.19 32.338 80 32.838 ;
        RECT 79.19 33.113 80 33.613 ;
        RECT 79.19 33.888 80 34.388 ;
        RECT 79.19 34.663 80 35.163 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C2 ;
        RECT 78.15 25 80 27.5 ;
      LAYER C1 ;
        RECT 79.19 24.838 80 27.663 ;
      LAYER M2 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER M1 ;
        RECT 79.19 24.838 80 25.338 ;
        RECT 79.19 25.613 80 26.113 ;
        RECT 79.19 26.388 80 26.888 ;
        RECT 79.19 27.163 80 27.663 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C2 ;
        RECT 78.15 10 80 12.5 ;
      LAYER C1 ;
        RECT 79.19 9.838 80 12.663 ;
      LAYER M2 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER M1 ;
        RECT 79.19 9.838 80 10.338 ;
        RECT 79.19 10.613 80 11.113 ;
        RECT 79.19 11.388 80 11.888 ;
        RECT 79.19 12.163 80 12.663 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSSX
  PIN VDDX
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddx VDDX!" ;
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C2 ;
        RECT 78.15 36.25 80 38.75 ;
      LAYER C1 ;
        RECT 79.19 36.088 80 38.913 ;
      LAYER M2 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
      LAYER M1 ;
        RECT 79.19 36.088 80 36.588 ;
        RECT 79.19 36.863 80 37.363 ;
        RECT 79.19 37.638 80 38.138 ;
        RECT 79.19 38.413 80 38.913 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C2 ;
        RECT 78.15 28.75 80 31.25 ;
      LAYER C1 ;
        RECT 79.19 28.588 80 31.413 ;
      LAYER M2 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
      LAYER M1 ;
        RECT 79.19 28.588 80 29.088 ;
        RECT 79.19 29.363 80 29.863 ;
        RECT 79.19 30.138 80 30.638 ;
        RECT 79.19 30.913 80 31.413 ;
    END
    PORT
      CLASS CORE ;
      LAYER C3 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C2 ;
        RECT 78.15 21.25 80 23.75 ;
      LAYER C1 ;
        RECT 79.19 21.088 80 23.913 ;
      LAYER M2 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
      LAYER M1 ;
        RECT 79.19 21.088 80 21.588 ;
        RECT 79.19 21.863 80 22.363 ;
        RECT 79.19 22.638 80 23.138 ;
        RECT 79.19 23.413 80 23.913 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C2 ;
        RECT 78.15 43.75 80 46.25 ;
      LAYER C1 ;
        RECT 79.19 43.588 80 46.413 ;
      LAYER M2 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER M1 ;
        RECT 79.19 43.588 80 44.088 ;
        RECT 79.19 44.363 80 44.863 ;
        RECT 79.19 45.138 80 45.638 ;
        RECT 79.19 45.913 80 46.413 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C2 ;
        RECT 78.15 13.75 80 16.25 ;
      LAYER C1 ;
        RECT 79.19 13.588 80 16.413 ;
      LAYER M2 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER M1 ;
        RECT 79.19 13.588 80 14.088 ;
        RECT 79.19 14.363 80 14.863 ;
        RECT 79.19 15.138 80 15.638 ;
        RECT 79.19 15.913 80 16.413 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
  END VDDX
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSSX_RVT_H

MACRO RIIO_EG1D80V_VSS_HVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS_HVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSS_HVT_H

MACRO RIIO_EG1D80V_VSS_RVT_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSS_RVT_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
    PORT
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSS_RVT_H

MACRO RIIO_EG1D80V_VSUP_CORE_GND_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_GND_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VSUP
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_CORE_GND_H

MACRO RIIO_EG1D80V_VSUP_CORE_PWR_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_PWR_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VSUP
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_CORE_PWR_H

MACRO RIIO_EG1D80V_VSUP_CORE_SIG_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_CORE_SIG_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.633 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1122.47 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 610.45 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 610.4525 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1151.7 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 770.45 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 454.315 LAYER IA ;
    ANTENNAPARTIALMETALAREA 397.03 LAYER IB ;
    ANTENNAPARTIALMETALAREA 4.554 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 2.392896 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 1.792 LAYER AY ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 26.515456 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 62.9856 LAYER YX ;
    ANTENNAPARTIALCUTAREA 40.310784 LAYER XA ;
    ANTENNAPARTIALCUTAREA 1.92 LAYER V1 ;
    ANTENNADIFFAREA 133.0532 LAYER C4 ;
    ANTENNADIFFAREA 133.0532 LAYER C3 ;
    ANTENNADIFFAREA 133.0532 LAYER C5 ;
    ANTENNADIFFAREA 133.0532 LAYER C6 ;
    ANTENNADIFFAREA 133.0532 LAYER IA ;
    ANTENNADIFFAREA 133.0532 LAYER IB ;
    ANTENNADIFFAREA 133.0532 LAYER C2 ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
        RECT 79.19 54.35 80 57.35 ;
    END
  END VSUP
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_CORE_SIG_H

MACRO RIIO_EG1D80V_VSUP_IO_GND_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_GND_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VSUP
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_IO_GND_H

MACRO RIIO_EG1D80V_VSUP_IO_PWR_H
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_PWR_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER IB ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER IA ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C6 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C5 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C4 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C3 ;
        RECT 0 49.35 1.85 52.95 ;
      LAYER C2 ;
        RECT 0 49.35 1.85 52.95 ;
    END
    PORT
      LAYER IB ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER IA ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C6 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C5 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C4 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C3 ;
        RECT 0 44.65 1.85 48.25 ;
      LAYER C2 ;
        RECT 0 44.65 1.85 48.25 ;
    END
    PORT
      LAYER IB ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER IA ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C6 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C5 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C4 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C3 ;
        RECT 0 39.95 1.85 43.55 ;
      LAYER C2 ;
        RECT 0 39.95 1.85 43.55 ;
    END
    PORT
      LAYER IB ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER IA ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C6 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C5 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C4 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C3 ;
        RECT 0 35.25 1.85 38.85 ;
      LAYER C2 ;
        RECT 0 35.25 1.85 38.85 ;
    END
    PORT
      LAYER IB ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER IA ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C6 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C5 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C4 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C3 ;
        RECT 0 30.55 1.85 34.15 ;
      LAYER C2 ;
        RECT 0 30.55 1.85 34.15 ;
    END
    PORT
      LAYER IB ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER IA ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C6 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C5 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C4 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C3 ;
        RECT 0 25.85 1.85 29.45 ;
      LAYER C2 ;
        RECT 0 25.85 1.85 29.45 ;
    END
    PORT
      LAYER IB ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER IA ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C6 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C5 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C4 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C3 ;
        RECT 0 21.15 1.85 24.75 ;
      LAYER C2 ;
        RECT 0 21.15 1.85 24.75 ;
    END
    PORT
      LAYER IB ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER IA ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C6 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C5 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C4 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C3 ;
        RECT 0 16.45 1.85 20.05 ;
      LAYER C2 ;
        RECT 0 16.45 1.85 20.05 ;
    END
    PORT
      LAYER IB ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER IA ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C6 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C5 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C4 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C3 ;
        RECT 0 11.75 1.85 15.35 ;
      LAYER C2 ;
        RECT 0 11.75 1.85 15.35 ;
    END
    PORT
      LAYER IB ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER IA ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C6 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C5 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C4 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C3 ;
        RECT 0 7.05 1.85 10.65 ;
      LAYER C2 ;
        RECT 0 7.05 1.85 10.65 ;
    END
    PORT
      LAYER IB ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
    END
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C2 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 54.35 80 57.35 ;
      LAYER M2 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M1 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER IA ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C6 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C5 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C4 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C3 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C2 ;
        RECT 78.15 49.65 80 52.65 ;
      LAYER C1 ;
        RECT 79.19 49.65 80 52.65 ;
      LAYER M2 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
      LAYER M1 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER IA ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C6 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C5 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C4 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C3 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C2 ;
        RECT 78.15 44.95 80 47.95 ;
      LAYER C1 ;
        RECT 79.19 44.95 80 47.95 ;
      LAYER M2 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
      LAYER M1 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER IA ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C6 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C5 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C4 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C3 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C2 ;
        RECT 78.15 40.25 80 43.25 ;
      LAYER C1 ;
        RECT 79.19 40.25 80 43.25 ;
      LAYER M2 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
      LAYER M1 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER IA ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C6 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C5 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C4 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C3 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C2 ;
        RECT 78.15 35.55 80 38.55 ;
      LAYER C1 ;
        RECT 79.19 35.55 80 38.55 ;
      LAYER M2 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
      LAYER M1 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER IA ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C6 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C5 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C4 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C3 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C2 ;
        RECT 78.15 30.85 80 33.85 ;
      LAYER C1 ;
        RECT 79.19 30.85 80 33.85 ;
      LAYER M2 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
      LAYER M1 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER IA ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C6 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C5 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C4 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C3 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C2 ;
        RECT 78.15 26.15 80 29.15 ;
      LAYER C1 ;
        RECT 79.19 26.15 80 29.15 ;
      LAYER M2 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
      LAYER M1 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER IA ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C6 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C5 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C4 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C3 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C2 ;
        RECT 78.15 21.45 80 24.45 ;
      LAYER C1 ;
        RECT 79.19 21.45 80 24.45 ;
      LAYER M2 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
      LAYER M1 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER IA ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C6 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C5 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C4 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C3 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C2 ;
        RECT 78.15 16.75 80 19.75 ;
      LAYER C1 ;
        RECT 79.19 16.75 80 19.75 ;
      LAYER M2 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
      LAYER M1 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER IA ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C6 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C5 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C4 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C3 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C2 ;
        RECT 78.15 12.05 80 15.05 ;
      LAYER C1 ;
        RECT 79.19 12.05 80 15.05 ;
      LAYER M2 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
      LAYER M1 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER IA ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C6 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C5 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C4 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C3 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C2 ;
        RECT 78.15 7.35 80 10.35 ;
      LAYER C1 ;
        RECT 79.19 7.35 80 10.35 ;
      LAYER M2 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
      LAYER M1 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
    END
  END VSUP
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_IO_PWR_H

MACRO RIIO_EG1D80V_VSUP_IO_SIG_H
  CLASS PAD INOUT ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_EG1D80V_VSUP_IO_SIG_H 0 0 ;
  SIZE 80 BY 60 ;
  SYMMETRY X Y ;
  SITE IO_EW_site ;
  PIN VSUP
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.633 LAYER C1 ;
    ANTENNAPARTIALMETALAREA 0.0495 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1151.7 LAYER C2 ;
    ANTENNAPARTIALMETALAREA 747.95 LAYER C3 ;
    ANTENNAPARTIALMETALAREA 611.5625 LAYER C4 ;
    ANTENNAPARTIALMETALAREA 1151.7 LAYER C5 ;
    ANTENNAPARTIALMETALAREA 770.45 LAYER C6 ;
    ANTENNAPARTIALMETALAREA 461.53 LAYER IA ;
    ANTENNAPARTIALMETALAREA 398.14 LAYER IB ;
    ANTENNAPARTIALMETALAREA 4.554 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 2.392896 LAYER A1 ;
    ANTENNAPARTIALCUTAREA 1.792 LAYER AY ;
    ANTENNAPARTIALCUTAREA 26.515456 LAYER A2 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A3 ;
    ANTENNAPARTIALCUTAREA 23.534016 LAYER A4 ;
    ANTENNAPARTIALCUTAREA 26.515456 LAYER A5 ;
    ANTENNAPARTIALCUTAREA 62.9856 LAYER YX ;
    ANTENNAPARTIALCUTAREA 40.310784 LAYER XA ;
    ANTENNAPARTIALCUTAREA 1.92 LAYER V1 ;
    ANTENNADIFFAREA 148.5876 LAYER C4 ;
    ANTENNADIFFAREA 148.5876 LAYER C3 ;
    ANTENNADIFFAREA 148.5876 LAYER C5 ;
    ANTENNADIFFAREA 148.5876 LAYER C6 ;
    ANTENNADIFFAREA 148.5876 LAYER IA ;
    ANTENNADIFFAREA 148.5876 LAYER IB ;
    ANTENNADIFFAREA 148.5876 LAYER C2 ;
    PORT
      LAYER IB ;
        RECT 21.75 2.35 25.35 57.65 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER IA ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C6 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C5 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C4 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C3 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
      LAYER C2 ;
        RECT 0 2.35 1.85 5.95 ;
        RECT 0 7.05 1.85 10.65 ;
        RECT 0 11.75 1.85 15.35 ;
        RECT 0 16.45 1.85 20.05 ;
        RECT 0 21.15 1.85 24.75 ;
        RECT 0 25.85 1.85 29.45 ;
        RECT 0 30.55 1.85 34.15 ;
        RECT 0 35.25 1.85 38.85 ;
        RECT 0 39.95 1.85 43.55 ;
        RECT 0 44.65 1.85 48.25 ;
        RECT 0 49.35 1.85 52.95 ;
        RECT 0 54.05 1.85 57.65 ;
    END
    PORT
      CLASS CORE ;
      LAYER IB ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER IA ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C6 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C5 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C4 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C3 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER M1 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER M2 ;
        RECT 79.19 2.35 80 2.85 ;
        RECT 79.19 3.125 80 3.625 ;
        RECT 79.19 3.9 80 4.4 ;
        RECT 79.19 4.675 80 5.175 ;
        RECT 79.19 5.45 80 5.95 ;
        RECT 79.19 7.05 80 7.55 ;
        RECT 79.19 7.825 80 8.325 ;
        RECT 79.19 8.6 80 9.1 ;
        RECT 79.19 9.375 80 9.875 ;
        RECT 79.19 10.15 80 10.65 ;
        RECT 79.19 11.75 80 12.25 ;
        RECT 79.19 12.525 80 13.025 ;
        RECT 79.19 13.3 80 13.8 ;
        RECT 79.19 14.075 80 14.575 ;
        RECT 79.19 14.85 80 15.35 ;
        RECT 79.19 16.45 80 16.95 ;
        RECT 79.19 17.225 80 17.725 ;
        RECT 79.19 18 80 18.5 ;
        RECT 79.19 18.775 80 19.275 ;
        RECT 79.19 19.55 80 20.05 ;
        RECT 79.19 21.15 80 21.65 ;
        RECT 79.19 21.925 80 22.425 ;
        RECT 79.19 22.7 80 23.2 ;
        RECT 79.19 23.475 80 23.975 ;
        RECT 79.19 24.25 80 24.75 ;
        RECT 79.19 25.85 80 26.35 ;
        RECT 79.19 26.625 80 27.125 ;
        RECT 79.19 27.4 80 27.9 ;
        RECT 79.19 28.175 80 28.675 ;
        RECT 79.19 28.95 80 29.45 ;
        RECT 79.19 30.55 80 31.05 ;
        RECT 79.19 31.325 80 31.825 ;
        RECT 79.19 32.1 80 32.6 ;
        RECT 79.19 32.875 80 33.375 ;
        RECT 79.19 33.65 80 34.15 ;
        RECT 79.19 35.25 80 35.75 ;
        RECT 79.19 36.025 80 36.525 ;
        RECT 79.19 36.8 80 37.3 ;
        RECT 79.19 37.575 80 38.075 ;
        RECT 79.19 38.35 80 38.85 ;
        RECT 79.19 39.95 80 40.45 ;
        RECT 79.19 40.725 80 41.225 ;
        RECT 79.19 41.5 80 42 ;
        RECT 79.19 42.275 80 42.775 ;
        RECT 79.19 43.05 80 43.55 ;
        RECT 79.19 44.65 80 45.15 ;
        RECT 79.19 45.425 80 45.925 ;
        RECT 79.19 46.2 80 46.7 ;
        RECT 79.19 46.975 80 47.475 ;
        RECT 79.19 47.75 80 48.25 ;
        RECT 79.19 49.35 80 49.85 ;
        RECT 79.19 50.125 80 50.625 ;
        RECT 79.19 50.9 80 51.4 ;
        RECT 79.19 51.675 80 52.175 ;
        RECT 79.19 52.45 80 52.95 ;
        RECT 79.19 54.05 80 54.55 ;
        RECT 79.19 54.825 80 55.325 ;
        RECT 79.19 55.6 80 56.1 ;
        RECT 79.19 56.375 80 56.875 ;
        RECT 79.19 57.15 80 57.65 ;
      LAYER C2 ;
        RECT 78.15 2.65 80 5.65 ;
        RECT 78.15 7.35 80 10.35 ;
        RECT 78.15 12.05 80 15.05 ;
        RECT 78.15 16.75 80 19.75 ;
        RECT 78.15 21.45 80 24.45 ;
        RECT 78.15 26.15 80 29.15 ;
        RECT 78.15 30.85 80 33.85 ;
        RECT 78.15 35.55 80 38.55 ;
        RECT 78.15 40.25 80 43.25 ;
        RECT 78.15 44.95 80 47.95 ;
        RECT 78.15 49.65 80 52.65 ;
        RECT 78.15 54.35 80 57.35 ;
      LAYER C1 ;
        RECT 79.19 2.65 80 5.65 ;
        RECT 79.19 7.35 80 10.35 ;
        RECT 79.19 12.05 80 15.05 ;
        RECT 79.19 16.75 80 19.75 ;
        RECT 79.19 21.45 80 24.45 ;
        RECT 79.19 26.15 80 29.15 ;
        RECT 79.19 30.85 80 33.85 ;
        RECT 79.19 35.55 80 38.55 ;
        RECT 79.19 40.25 80 43.25 ;
        RECT 79.19 44.95 80 47.95 ;
        RECT 79.19 49.65 80 52.65 ;
        RECT 79.19 54.35 80 57.35 ;
    END
  END VSUP
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER IB ;
        RECT 59.35 0 62.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 73.45 0 77.05 60 ;
    END
  END VSS
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddio VDDIO!" ;
    PORT
      LAYER IB ;
        RECT 7.65 0 11.25 60 ;
    END
    PORT
      LAYER IB ;
        RECT 12.35 0 15.95 60 ;
    END
    PORT
      LAYER IB ;
        RECT 31.15 0 34.75 60 ;
    END
    PORT
      LAYER IB ;
        RECT 35.85 0 39.45 60 ;
    END
    PORT
      LAYER IB ;
        RECT 49.95 0 53.55 60 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vssio VSSIO!" ;
    PORT
      LAYER IB ;
        RECT 3.67 0 6.55 60 ;
    END
    PORT
      LAYER IB ;
        RECT 17.05 0 20.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 26.45 0 30.05 60 ;
    END
    PORT
      LAYER IB ;
        RECT 40.55 0 44.15 60 ;
    END
    PORT
      LAYER IB ;
        RECT 45.25 0 48.85 60 ;
    END
    PORT
      LAYER IB ;
        RECT 54.65 0 58.25 60 ;
    END
  END VSSIO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER IB ;
        RECT 64.05 0 67.65 60 ;
    END
    PORT
      LAYER IB ;
        RECT 68.75 0 72.35 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 60 ;
    LAYER M1 ;
      RECT 0 0 80 60 ;
    LAYER V1 ;
      RECT 0 0 80 60 ;
    LAYER M2 ;
      RECT 0 0 80 60 ;
    LAYER A1 ;
      RECT 0 0 80 60 ;
    LAYER C2 ;
      RECT 0 0 80 60 ;
    LAYER IA ;
      RECT 0 0 80 60 ;
    LAYER XA ;
      RECT 0 0 80 60 ;
    LAYER YX ;
      RECT 0 0 80 60 ;
    LAYER IB ;
      RECT 0 0 80 60 ;
    LAYER CB ;
      RECT 0 0 80 60 ;
    LAYER AY ;
      RECT 0 0 80 60 ;
    LAYER C1 ;
      RECT 0 0 80 60 ;
    LAYER C5 ;
      RECT 0 0 80 60 ;
    LAYER C4 ;
      RECT 0 0 80 60 ;
    LAYER C3 ;
      RECT 0 0 80 60 ;
    LAYER A5 ;
      RECT 0 0 80 60 ;
    LAYER A4 ;
      RECT 0 0 80 60 ;
    LAYER A3 ;
      RECT 0 0 80 60 ;
    LAYER A2 ;
      RECT 0 0 80 60 ;
    LAYER C6 ;
      RECT 0 0 80 60 ;
  END
END RIIO_EG1D80V_VSUP_IO_SIG_H





















MACRO RIIO_BOND20x10_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND20x10_INNER_GND 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 10.01 0 29.99 10 ;
      LAYER IB ;
        RECT 15 0 25 10 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER IA ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 10 5 29.99 10 ;
      RECT 10.01 0 30 5 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER XA ;
      RECT 0 0 40 10 ;
    LAYER YX ;
      RECT 0 0 40 10 ;
    LAYER IB ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A5 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
    LAYER C6 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND20x10_INNER_GND

MACRO RIIO_BOND20x10_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND20x10_INNER_PWR 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 10 0 30 10 ;
      LAYER IB ;
        RECT 15 0 25 10 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER IA ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 10 0 30 10 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER XA ;
      RECT 0 0 40 10 ;
    LAYER YX ;
      RECT 0 0 40 10 ;
    LAYER IB ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A5 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
    LAYER C6 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND20x10_INNER_PWR

MACRO RIIO_BOND20x10_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND20x10_INNER_SIG 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 206.8788 LAYER IB ;
    ANTENNAPARTIALCUTAREA 43.74 LAYER VV ;
    PORT
      LAYER IB ;
        RECT 15 0 25 10 ;
      LAYER LB ;
        RECT 10 0 30 10 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER IA ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 10 0 30 10 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER XA ;
      RECT 0 0 40 10 ;
    LAYER YX ;
      RECT 0 0 40 10 ;
    LAYER IB ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A5 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
    LAYER C6 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND20x10_INNER_SIG

MACRO RIIO_BOND60_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_INNER_GND 0 0 ;
  SIZE 60 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 10 0 50 70 ;
      LAYER IB ;
        RECT 10 69 50 70 ;
      LAYER IA ;
        RECT 10 69 50 70 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER IA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER XA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER YX ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER IB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A5 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C6 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  50 60  50 70  10 70  10 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_INNER_GND

MACRO RIIO_BOND60_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_INNER_PWR 0 0 ;
  SIZE 60 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 10 0 50 70 ;
      LAYER IB ;
        RECT 10 69 50 70 ;
      LAYER IA ;
        RECT 10 69 50 70 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER IA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER XA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER YX ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER IB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A5 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C6 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  50 60  50 70  10 70  10 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_INNER_PWR

MACRO RIIO_BOND60_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_INNER_SIG 0 0 ;
  SIZE 60 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2497.68 LAYER IA ;
    ANTENNAPARTIALMETALAREA 2950.18 LAYER IB ;
    ANTENNAPARTIALCUTAREA 379.173312 LAYER XA ;
    ANTENNAPARTIALCUTAREA 408.24 LAYER VV ;
    PORT
      LAYER IA ;
        RECT 10 69 50 70 ;
      LAYER IB ;
        RECT 10 69 50 70 ;
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 10 0 50 70 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER IA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER XA ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER YX ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER IB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A5 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER C6 ;
      RECT 10 0 50 70 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  50 60  50 70  10 70  10 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_INNER_SIG

MACRO RIIO_BOND60_OUTER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_OUTER_GND 0 0 ;
  SIZE 60 BY 140 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 12.5 0 47.5 140 ;
      LAYER IB ;
        RECT 12.5 139 47.5 140 ;
      LAYER IA ;
        RECT 12.5 139 47.5 140 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER IA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER XA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER YX ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER IB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A5 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C6 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  47.5 60  47.5 140  12.5 140  12.5 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_OUTER_GND

MACRO RIIO_BOND60_OUTER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_OUTER_PWR 0 0 ;
  SIZE 60 BY 140 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 12.5 0 47.5 140 ;
      LAYER IB ;
        RECT 12.5 139 47.5 140 ;
      LAYER IA ;
        RECT 12.5 139 47.5 140 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER IA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER XA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER YX ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER IB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A5 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C6 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  47.5 60  47.5 140  12.5 140  12.5 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_OUTER_PWR

MACRO RIIO_BOND60_OUTER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_OUTER_SIG 0 0 ;
  SIZE 60 BY 140 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3588.5016 LAYER IA ;
    ANTENNAPARTIALMETALAREA 4731.2304 LAYER IB ;
    ANTENNAPARTIALCUTAREA 559.312128 LAYER XA ;
    ANTENNAPARTIALCUTAREA 903.96 LAYER VV ;
    PORT
      LAYER IA ;
        RECT 12.5 139 47.5 140 ;
      LAYER IB ;
        RECT 12.5 139 47.5 140 ;
      LAYER LB ;
        RECT 0 0 60 60 ;
        RECT 12.5 0 47.5 140 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER IA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER XA ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER YX ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER IB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A5 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER C6 ;
      RECT 12.5 0 47.5 140 ;
      RECT 0 0 60 60 ;
    LAYER OVERLAP ;
      POLYGON  60 60  47.5 60  47.5 140  12.5 140  12.5 60  0 60  0 0  60 0 ;
  END
END RIIO_BOND60_OUTER_SIG

MACRO RIIO_BOND60_PLAIN_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_PLAIN_GND 0 0 ;
  SIZE 60 BY 60 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 0 0 60 60 ;
    LAYER IA ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 0 0 60 60 ;
    LAYER XA ;
      RECT 0 0 60 60 ;
    LAYER YX ;
      RECT 0 0 60 60 ;
    LAYER IB ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 0 0 60 60 ;
    LAYER A5 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 0 0 60 60 ;
    LAYER C6 ;
      RECT 0 0 60 60 ;
  END
END RIIO_BOND60_PLAIN_GND

MACRO RIIO_BOND60_PLAIN_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_PLAIN_PWR 0 0 ;
  SIZE 60 BY 60 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 0 0 60 60 ;
    LAYER IA ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 0 0 60 60 ;
    LAYER XA ;
      RECT 0 0 60 60 ;
    LAYER YX ;
      RECT 0 0 60 60 ;
    LAYER IB ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 0 0 60 60 ;
    LAYER A5 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 0 0 60 60 ;
    LAYER C6 ;
      RECT 0 0 60 60 ;
  END
END RIIO_BOND60_PLAIN_PWR

MACRO RIIO_BOND60_PLAIN_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60_PLAIN_SIG 0 0 ;
  SIZE 60 BY 60 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 60 60 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 60 60 ;
    LAYER M1 ;
      RECT 0 0 60 60 ;
    LAYER V1 ;
      RECT 0 0 60 60 ;
    LAYER M2 ;
      RECT 0 0 60 60 ;
    LAYER A1 ;
      RECT 0 0 60 60 ;
    LAYER C2 ;
      RECT 0 0 60 60 ;
    LAYER IA ;
      RECT 0 0 60 60 ;
    LAYER LB ;
      RECT 0 0 60 60 ;
    LAYER VV ;
      RECT 0 0 60 60 ;
    LAYER XA ;
      RECT 0 0 60 60 ;
    LAYER YX ;
      RECT 0 0 60 60 ;
    LAYER IB ;
      RECT 0 0 60 60 ;
    LAYER CB ;
      RECT 0 0 60 60 ;
    LAYER AY ;
      RECT 0 0 60 60 ;
    LAYER C1 ;
      RECT 0 0 60 60 ;
    LAYER C5 ;
      RECT 0 0 60 60 ;
    LAYER C4 ;
      RECT 0 0 60 60 ;
    LAYER C3 ;
      RECT 0 0 60 60 ;
    LAYER A5 ;
      RECT 0 0 60 60 ;
    LAYER A4 ;
      RECT 0 0 60 60 ;
    LAYER A3 ;
      RECT 0 0 60 60 ;
    LAYER A2 ;
      RECT 0 0 60 60 ;
    LAYER C6 ;
      RECT 0 0 60 60 ;
  END
END RIIO_BOND60_PLAIN_SIG

MACRO RIIO_BOND60x90_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_GND 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
      LAYER IB ;
        RECT 10 99 50 100 ;
      LAYER IA ;
        RECT 10 99 50 100 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_GND

MACRO RIIO_BOND60x90_INNER_GND_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_GND_CESD 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
      LAYER IB ;
        RECT 10 99 50 100 ;
      LAYER IA ;
        RECT 10 99 50 100 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_GND_CESD

MACRO RIIO_BOND60x90_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_PWR 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
      LAYER IB ;
        RECT 10 99 50 100 ;
      LAYER IA ;
        RECT 10 99 50 100 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_PWR

MACRO RIIO_BOND60x90_INNER_PWR_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_PWR_CESD 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
      LAYER IB ;
        RECT 10 99 50 100 ;
      LAYER IA ;
        RECT 10 99 50 100 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_PWR_CESD

MACRO RIIO_BOND60x90_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_SIG 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3797.68 LAYER IA ;
    ANTENNAPARTIALMETALAREA 4370.18 LAYER IB ;
    ANTENNAPARTIALCUTAREA 564.350976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 495.72 LAYER VV ;
    PORT
      LAYER IA ;
        RECT 10 99 50 100 ;
      LAYER IB ;
        RECT 10 99 50 100 ;
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_SIG

MACRO RIIO_BOND60x90_INNER_SIG_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_INNER_SIG_CESD 0 0 ;
  SIZE 60 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3797.68 LAYER IA ;
    ANTENNAPARTIALMETALAREA 4370.18 LAYER IB ;
    ANTENNAPARTIALCUTAREA 564.350976 LAYER XA ;
    ANTENNAPARTIALCUTAREA 495.72 LAYER VV ;
    PORT
      LAYER IA ;
        RECT 10 99 50 100 ;
      LAYER IB ;
        RECT 10 99 50 100 ;
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 10 0 50 100 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 10 0 50 100 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  50 90  50 100  10 100  10 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_INNER_SIG_CESD

MACRO RIIO_BOND60x90_OUTER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_GND 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
      LAYER IB ;
        RECT 12.5 199 47.5 200 ;
      LAYER IA ;
        RECT 12.5 199 47.5 200 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_GND

MACRO RIIO_BOND60x90_OUTER_GND_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_GND_CESD 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
      LAYER IB ;
        RECT 12.5 199 47.5 200 ;
      LAYER IA ;
        RECT 12.5 199 47.5 200 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_GND_CESD

MACRO RIIO_BOND60x90_OUTER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_PWR 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
      LAYER IB ;
        RECT 12.5 199 47.5 200 ;
      LAYER IA ;
        RECT 12.5 199 47.5 200 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_PWR

MACRO RIIO_BOND60x90_OUTER_PWR_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_PWR_CESD 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
      LAYER IB ;
        RECT 12.5 199 47.5 200 ;
      LAYER IA ;
        RECT 12.5 199 47.5 200 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_PWR_CESD

MACRO RIIO_BOND60x90_OUTER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_SIG 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5221.2668 LAYER IA ;
    ANTENNAPARTIALMETALAREA 6933.5668 LAYER IB ;
    ANTENNAPARTIALCUTAREA 823.851648 LAYER XA ;
    ANTENNAPARTIALCUTAREA 1210.14 LAYER VV ;
    PORT
      LAYER IA ;
        RECT 12.5 199 47.5 200 ;
      LAYER IB ;
        RECT 12.5 199 47.5 200 ;
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_SIG

MACRO RIIO_BOND60x90_OUTER_SIG_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_OUTER_SIG_CESD 0 0 ;
  SIZE 60 BY 200 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5221.2668 LAYER IA ;
    ANTENNAPARTIALMETALAREA 6933.5668 LAYER IB ;
    ANTENNAPARTIALCUTAREA 823.851648 LAYER XA ;
    ANTENNAPARTIALCUTAREA 1210.14 LAYER VV ;
    PORT
      LAYER IA ;
        RECT 12.5 199 47.5 200 ;
      LAYER IB ;
        RECT 12.5 199 47.5 200 ;
      LAYER LB ;
        RECT 0 0 60 90 ;
        RECT 12.5 0 47.5 200 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 12.5 0 47.5 200 ;
      RECT 0 0 60 90 ;
    LAYER OVERLAP ;
      POLYGON  60 90  47.5 90  47.5 200  12.5 200  12.5 90  0 90  0 0  60 0 ;
  END
END RIIO_BOND60x90_OUTER_SIG_CESD

MACRO RIIO_BOND60x90_PLAIN_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_GND 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_GND

MACRO RIIO_BOND60x90_PLAIN_GND_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_GND_CESD 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_GND_CESD

MACRO RIIO_BOND60x90_PLAIN_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_PWR 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_PWR

MACRO RIIO_BOND60x90_PLAIN_PWR_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_PWR_CESD 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_PWR_CESD

MACRO RIIO_BOND60x90_PLAIN_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_SIG 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_SIG

MACRO RIIO_BOND60x90_PLAIN_SIG_CESD
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND60x90_PLAIN_SIG_CESD 0 0 ;
  SIZE 60 BY 90 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 60 90 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 60 90 ;
    LAYER M1 ;
      RECT 0 0 60 90 ;
    LAYER V1 ;
      RECT 0 0 60 90 ;
    LAYER M2 ;
      RECT 0 0 60 90 ;
    LAYER A1 ;
      RECT 0 0 60 90 ;
    LAYER C2 ;
      RECT 0 0 60 90 ;
    LAYER IA ;
      RECT 0 0 60 90 ;
    LAYER LB ;
      RECT 0 0 60 90 ;
    LAYER VV ;
      RECT 0 0 60 90 ;
    LAYER XA ;
      RECT 0 0 60 90 ;
    LAYER YX ;
      RECT 0 0 60 90 ;
    LAYER IB ;
      RECT 0 0 60 90 ;
    LAYER CB ;
      RECT 0 0 60 90 ;
    LAYER AY ;
      RECT 0 0 60 90 ;
    LAYER C1 ;
      RECT 0 0 60 90 ;
    LAYER C5 ;
      RECT 0 0 60 90 ;
    LAYER C4 ;
      RECT 0 0 60 90 ;
    LAYER C3 ;
      RECT 0 0 60 90 ;
    LAYER A5 ;
      RECT 0 0 60 90 ;
    LAYER A4 ;
      RECT 0 0 60 90 ;
    LAYER A3 ;
      RECT 0 0 60 90 ;
    LAYER A2 ;
      RECT 0 0 60 90 ;
    LAYER C6 ;
      RECT 0 0 60 90 ;
  END
END RIIO_BOND60x90_PLAIN_SIG_CESD

MACRO RIIO_BOND64_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_INNER_GND 0 0 ;
  SIZE 64 BY 72 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 12 0 52 72 ;
      LAYER IB ;
        RECT 12 71 52 72 ;
      LAYER IA ;
        RECT 12 71 52 72 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER IA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER XA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER YX ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER IB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A5 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C6 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 72  12 72  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_INNER_GND

MACRO RIIO_BOND64_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_INNER_PWR 0 0 ;
  SIZE 64 BY 72 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 12 0 52 72 ;
      LAYER IB ;
        RECT 12 71 52 72 ;
      LAYER IA ;
        RECT 12 71 52 72 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER IA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER XA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER YX ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER IB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A5 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C6 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 72  12 72  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_INNER_PWR

MACRO RIIO_BOND64_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_INNER_SIG 0 0 ;
  SIZE 64 BY 72 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2746.5 LAYER IA ;
    ANTENNAPARTIALMETALAREA 3083.5 LAYER IB ;
    ANTENNAPARTIALCUTAREA 436.490208 LAYER XA ;
    ANTENNAPARTIALCUTAREA 408.24 LAYER VV ;
    PORT
      LAYER IA ;
        RECT 12 71 52 72 ;
      LAYER IB ;
        RECT 12 71 52 72 ;
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 12 0 52 72 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER IA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER XA ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER YX ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER IB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A5 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER C6 ;
      RECT 12 0 52 72 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 72  12 72  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_INNER_SIG

MACRO RIIO_BOND64_OUTER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_OUTER_GND 0 0 ;
  SIZE 64 BY 144 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 11.998 0 52 144 ;
      LAYER IB ;
        RECT 12 143 52 144 ;
      LAYER IA ;
        RECT 12 143 52 144 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER IA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 11.998 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER XA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER YX ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER IB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A5 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C6 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 144  12 144  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_OUTER_GND

MACRO RIIO_BOND64_OUTER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_OUTER_PWR 0 0 ;
  SIZE 64 BY 144 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 11.998 0 52 144 ;
      LAYER IB ;
        RECT 12 143 52 144 ;
      LAYER IA ;
        RECT 12 143 52 144 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER IA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 11.998 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER XA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER YX ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER IB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A5 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C6 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 144  12 144  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_OUTER_PWR

MACRO RIIO_BOND64_OUTER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_OUTER_SIG 0 0 ;
  SIZE 64 BY 144 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4096.5 LAYER IA ;
    ANTENNAPARTIALMETALAREA 4841.5 LAYER IB ;
    ANTENNAPARTIALCUTAREA 630.485856 LAYER XA ;
    ANTENNAPARTIALCUTAREA 816.48 LAYER VV ;
    PORT
      LAYER IA ;
        RECT 12 143 52 144 ;
      LAYER IB ;
        RECT 12 143 52 144 ;
      LAYER LB ;
        RECT 0 0 64 64 ;
        RECT 11.998 0 52 144 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER IA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 11.998 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER XA ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER YX ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER IB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A5 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER C6 ;
      RECT 12 0 52 144 ;
      RECT 0 0 64 64 ;
    LAYER OVERLAP ;
      POLYGON  64 64  52 64  52 144  12 144  12 64  0 64  0 0  64 0 ;
  END
END RIIO_BOND64_OUTER_SIG

MACRO RIIO_BOND64_PLAIN_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_PLAIN_GND 0 0 ;
  SIZE 64 BY 64 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 0 0 64 64 ;
    LAYER IA ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 0 0 64 64 ;
    LAYER XA ;
      RECT 0 0 64 64 ;
    LAYER YX ;
      RECT 0 0 64 64 ;
    LAYER IB ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 0 0 64 64 ;
    LAYER A5 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 0 0 64 64 ;
    LAYER C6 ;
      RECT 0 0 64 64 ;
  END
END RIIO_BOND64_PLAIN_GND

MACRO RIIO_BOND64_PLAIN_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_PLAIN_PWR 0 0 ;
  SIZE 64 BY 64 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 0 0 64 64 ;
    LAYER IA ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 0 0 64 64 ;
    LAYER XA ;
      RECT 0 0 64 64 ;
    LAYER YX ;
      RECT 0 0 64 64 ;
    LAYER IB ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 0 0 64 64 ;
    LAYER A5 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 0 0 64 64 ;
    LAYER C6 ;
      RECT 0 0 64 64 ;
  END
END RIIO_BOND64_PLAIN_PWR

MACRO RIIO_BOND64_PLAIN_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND64_PLAIN_SIG 0 0 ;
  SIZE 64 BY 64 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 64 64 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 64 64 ;
    LAYER M1 ;
      RECT 0 0 64 64 ;
    LAYER V1 ;
      RECT 0 0 64 64 ;
    LAYER M2 ;
      RECT 0 0 64 64 ;
    LAYER A1 ;
      RECT 0 0 64 64 ;
    LAYER C2 ;
      RECT 0 0 64 64 ;
    LAYER IA ;
      RECT 0 0 64 64 ;
    LAYER LB ;
      RECT 0 0 64 64 ;
    LAYER VV ;
      RECT 0 0 64 64 ;
    LAYER XA ;
      RECT 0 0 64 64 ;
    LAYER YX ;
      RECT 0 0 64 64 ;
    LAYER IB ;
      RECT 0 0 64 64 ;
    LAYER CB ;
      RECT 0 0 64 64 ;
    LAYER AY ;
      RECT 0 0 64 64 ;
    LAYER C1 ;
      RECT 0 0 64 64 ;
    LAYER C5 ;
      RECT 0 0 64 64 ;
    LAYER C4 ;
      RECT 0 0 64 64 ;
    LAYER C3 ;
      RECT 0 0 64 64 ;
    LAYER A5 ;
      RECT 0 0 64 64 ;
    LAYER A4 ;
      RECT 0 0 64 64 ;
    LAYER A3 ;
      RECT 0 0 64 64 ;
    LAYER A2 ;
      RECT 0 0 64 64 ;
    LAYER C6 ;
      RECT 0 0 64 64 ;
  END
END RIIO_BOND64_PLAIN_SIG

MACRO RIIO_BOND70_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_INNER_GND 0 0 ;
  SIZE 70 BY 80 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 15 0 55 80 ;
      LAYER IB ;
        RECT 15 79 55 80 ;
      LAYER IA ;
        RECT 15 79 55 80 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER IA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER XA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER YX ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER IB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A5 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C6 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  55 70  55 80  15 80  15 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_INNER_GND

MACRO RIIO_BOND70_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_INNER_PWR 0 0 ;
  SIZE 70 BY 80 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 15 0 55 80 ;
      LAYER IB ;
        RECT 15 79 55 80 ;
      LAYER IA ;
        RECT 15 79 55 80 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER IA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER XA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER YX ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER IB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A5 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C6 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  55 70  55 80  15 80  15 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_INNER_PWR

MACRO RIIO_BOND70_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_INNER_SIG 0 0 ;
  SIZE 70 BY 80 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3447.68 LAYER IA ;
    ANTENNAPARTIALMETALAREA 3975.18 LAYER IB ;
    ANTENNAPARTIALCUTAREA 522.78048 LAYER XA ;
    ANTENNAPARTIALCUTAREA 466.56 LAYER VV ;
    PORT
      LAYER IA ;
        RECT 15 79 55 80 ;
      LAYER IB ;
        RECT 15 79 55 80 ;
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 15 0 55 80 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER IA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER XA ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER YX ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER IB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A5 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER C6 ;
      RECT 15 0 55 80 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  55 70  55 80  15 80  15 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_INNER_SIG

MACRO RIIO_BOND70_OUTER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_OUTER_GND 0 0 ;
  SIZE 70 BY 160 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 17.5 0 52.5 160 ;
      LAYER IB ;
        RECT 17.5 159 52.5 160 ;
      LAYER IA ;
        RECT 17.5 159 52.5 160 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER IA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER XA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER YX ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER IB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A5 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C6 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  52.5 70  52.5 160  17.5 160  17.5 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_OUTER_GND

MACRO RIIO_BOND70_OUTER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_OUTER_PWR 0 0 ;
  SIZE 70 BY 160 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 17.5 0 52.5 160 ;
      LAYER IB ;
        RECT 17.5 159 52.5 160 ;
      LAYER IA ;
        RECT 17.5 159 52.5 160 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER IA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER XA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER YX ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER IB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A5 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C6 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  52.5 70  52.5 160  17.5 160  17.5 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_OUTER_PWR

MACRO RIIO_BOND70_OUTER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_OUTER_SIG 0 0 ;
  SIZE 70 BY 160 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4288.88 LAYER IA ;
    ANTENNAPARTIALMETALAREA 6011.62 LAYER IB ;
    ANTENNAPARTIALCUTAREA 729.373248 LAYER XA ;
    ANTENNAPARTIALCUTAREA 1035.18 LAYER VV ;
    PORT
      LAYER IA ;
        RECT 17.5 159 52.5 160 ;
      LAYER IB ;
        RECT 17.5 159 52.5 160 ;
      LAYER LB ;
        RECT 0 0 70 70 ;
        RECT 17.5 0 52.5 160 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER IA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER XA ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER YX ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER IB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A5 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER C6 ;
      RECT 17.5 0 52.5 160 ;
      RECT 0 0 70 70 ;
    LAYER OVERLAP ;
      POLYGON  70 70  52.5 70  52.5 160  17.5 160  17.5 70  0 70  0 0  70 0 ;
  END
END RIIO_BOND70_OUTER_SIG

MACRO RIIO_BOND70_PLAIN_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_PLAIN_GND 0 0 ;
  SIZE 70 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 0 0 70 70 ;
    LAYER IA ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 0 0 70 70 ;
    LAYER XA ;
      RECT 0 0 70 70 ;
    LAYER YX ;
      RECT 0 0 70 70 ;
    LAYER IB ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 0 0 70 70 ;
    LAYER A5 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 0 0 70 70 ;
    LAYER C6 ;
      RECT 0 0 70 70 ;
  END
END RIIO_BOND70_PLAIN_GND

MACRO RIIO_BOND70_PLAIN_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_PLAIN_PWR 0 0 ;
  SIZE 70 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 0 0 70 70 ;
    LAYER IA ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 0 0 70 70 ;
    LAYER XA ;
      RECT 0 0 70 70 ;
    LAYER YX ;
      RECT 0 0 70 70 ;
    LAYER IB ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 0 0 70 70 ;
    LAYER A5 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 0 0 70 70 ;
    LAYER C6 ;
      RECT 0 0 70 70 ;
  END
END RIIO_BOND70_PLAIN_PWR

MACRO RIIO_BOND70_PLAIN_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND70_PLAIN_SIG 0 0 ;
  SIZE 70 BY 70 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 70 70 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 70 70 ;
    LAYER M1 ;
      RECT 0 0 70 70 ;
    LAYER V1 ;
      RECT 0 0 70 70 ;
    LAYER M2 ;
      RECT 0 0 70 70 ;
    LAYER A1 ;
      RECT 0 0 70 70 ;
    LAYER C2 ;
      RECT 0 0 70 70 ;
    LAYER IA ;
      RECT 0 0 70 70 ;
    LAYER LB ;
      RECT 0 0 70 70 ;
    LAYER VV ;
      RECT 0 0 70 70 ;
    LAYER XA ;
      RECT 0 0 70 70 ;
    LAYER YX ;
      RECT 0 0 70 70 ;
    LAYER IB ;
      RECT 0 0 70 70 ;
    LAYER CB ;
      RECT 0 0 70 70 ;
    LAYER AY ;
      RECT 0 0 70 70 ;
    LAYER C1 ;
      RECT 0 0 70 70 ;
    LAYER C5 ;
      RECT 0 0 70 70 ;
    LAYER C4 ;
      RECT 0 0 70 70 ;
    LAYER C3 ;
      RECT 0 0 70 70 ;
    LAYER A5 ;
      RECT 0 0 70 70 ;
    LAYER A4 ;
      RECT 0 0 70 70 ;
    LAYER A3 ;
      RECT 0 0 70 70 ;
    LAYER A2 ;
      RECT 0 0 70 70 ;
    LAYER C6 ;
      RECT 0 0 70 70 ;
  END
END RIIO_BOND70_PLAIN_SIG

MACRO RIIO_BOND80x100_INNER_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_INNER_GND 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT -20 -110 60 -10 ;
        RECT 0 -110 40 10 ;
      LAYER IB ;
        RECT 15 0 25 10 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER IA ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 0 -110 40 10 ;
      RECT -20 -110 60 -10 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER XA ;
      RECT 0 0 40 10 ;
    LAYER YX ;
      RECT 0 0 40 10 ;
    LAYER IB ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A5 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
    LAYER C6 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND80x100_INNER_GND

MACRO RIIO_BOND80x100_INNER_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_INNER_PWR 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT -20 -110 60 -10 ;
        RECT 0 -110 40 10 ;
      LAYER IB ;
        RECT 15 0 25 10 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER IA ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 0 -110 40 10 ;
      RECT -20 -110 60 -10 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER XA ;
      RECT 0 0 40 10 ;
    LAYER YX ;
      RECT 0 0 40 10 ;
    LAYER IB ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A5 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
    LAYER C6 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND80x100_INNER_PWR

MACRO RIIO_BOND80x100_INNER_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_INNER_SIG 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.2576 LAYER IB ;
    ANTENNAPARTIALCUTAREA 29.16 LAYER VV ;
    PORT
      LAYER IB ;
        RECT 15 0 25 10 ;
      LAYER LB ;
        RECT -20 -110 60 -10 ;
        RECT 0 -110 40 10 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 40 10 ;
    LAYER M1 ;
      RECT 0 0 40 10 ;
    LAYER V1 ;
      RECT 0 0 40 10 ;
    LAYER M2 ;
      RECT 0 0 40 10 ;
    LAYER A1 ;
      RECT 0 0 40 10 ;
    LAYER C2 ;
      RECT 0 0 40 10 ;
    LAYER IA ;
      RECT 0 0 40 10 ;
    LAYER LB ;
      RECT 0 -110 40 10 ;
      RECT -20 -110 60 -10 ;
    LAYER VV ;
      RECT 0 0 40 10 ;
    LAYER XA ;
      RECT 0 0 40 10 ;
    LAYER YX ;
      RECT 0 0 40 10 ;
    LAYER IB ;
      RECT 0 0 40 10 ;
    LAYER CB ;
      RECT 0 0 40 10 ;
    LAYER AY ;
      RECT 0 0 40 10 ;
    LAYER C1 ;
      RECT 0 0 40 10 ;
    LAYER C5 ;
      RECT 0 0 40 10 ;
    LAYER C4 ;
      RECT 0 0 40 10 ;
    LAYER C3 ;
      RECT 0 0 40 10 ;
    LAYER A5 ;
      RECT 0 0 40 10 ;
    LAYER A4 ;
      RECT 0 0 40 10 ;
    LAYER A3 ;
      RECT 0 0 40 10 ;
    LAYER A2 ;
      RECT 0 0 40 10 ;
    LAYER C6 ;
      RECT 0 0 40 10 ;
  END
END RIIO_BOND80x100_INNER_SIG

MACRO RIIO_BOND80x100_PLAIN_GND
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_PLAIN_GND 0 0 ;
  SIZE 80 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
        RECT 0 0 80 100 ;
    END
  END VSS
  OBS
    LAYER CA ;
      RECT 0 0 80 100 ;
    LAYER M1 ;
      RECT 0 0 80 100 ;
    LAYER V1 ;
      RECT 0 0 80 100 ;
    LAYER M2 ;
      RECT 0 0 80 100 ;
    LAYER A1 ;
      RECT 0 0 80 100 ;
    LAYER C2 ;
      RECT 0 0 80 100 ;
    LAYER IA ;
      RECT 0 0 80 100 ;
    LAYER LB ;
      RECT 0 0 80 100 ;
    LAYER VV ;
      RECT 0 0 80 100 ;
    LAYER XA ;
      RECT 0 0 80 100 ;
    LAYER YX ;
      RECT 0 0 80 100 ;
    LAYER IB ;
      RECT 0 0 80 100 ;
    LAYER CB ;
      RECT 0 0 80 100 ;
    LAYER AY ;
      RECT 0 0 80 100 ;
    LAYER C1 ;
      RECT 0 0 80 100 ;
    LAYER C5 ;
      RECT 0 0 80 100 ;
    LAYER C4 ;
      RECT 0 0 80 100 ;
    LAYER C3 ;
      RECT 0 0 80 100 ;
    LAYER A5 ;
      RECT 0 0 80 100 ;
    LAYER A4 ;
      RECT 0 0 80 100 ;
    LAYER A3 ;
      RECT 0 0 80 100 ;
    LAYER A2 ;
      RECT 0 0 80 100 ;
    LAYER C6 ;
      RECT 0 0 80 100 ;
  END
END RIIO_BOND80x100_PLAIN_GND

MACRO RIIO_BOND80x100_PLAIN_PWR
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_PLAIN_PWR 0 0 ;
  SIZE 80 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
        RECT 0 0 80 100 ;
    END
  END VDD
  OBS
    LAYER CA ;
      RECT 0 0 80 100 ;
    LAYER M1 ;
      RECT 0 0 80 100 ;
    LAYER V1 ;
      RECT 0 0 80 100 ;
    LAYER M2 ;
      RECT 0 0 80 100 ;
    LAYER A1 ;
      RECT 0 0 80 100 ;
    LAYER C2 ;
      RECT 0 0 80 100 ;
    LAYER IA ;
      RECT 0 0 80 100 ;
    LAYER LB ;
      RECT 0 0 80 100 ;
    LAYER VV ;
      RECT 0 0 80 100 ;
    LAYER XA ;
      RECT 0 0 80 100 ;
    LAYER YX ;
      RECT 0 0 80 100 ;
    LAYER IB ;
      RECT 0 0 80 100 ;
    LAYER CB ;
      RECT 0 0 80 100 ;
    LAYER AY ;
      RECT 0 0 80 100 ;
    LAYER C1 ;
      RECT 0 0 80 100 ;
    LAYER C5 ;
      RECT 0 0 80 100 ;
    LAYER C4 ;
      RECT 0 0 80 100 ;
    LAYER C3 ;
      RECT 0 0 80 100 ;
    LAYER A5 ;
      RECT 0 0 80 100 ;
    LAYER A4 ;
      RECT 0 0 80 100 ;
    LAYER A3 ;
      RECT 0 0 80 100 ;
    LAYER A2 ;
      RECT 0 0 80 100 ;
    LAYER C6 ;
      RECT 0 0 80 100 ;
  END
END RIIO_BOND80x100_PLAIN_PWR

MACRO RIIO_BOND80x100_PLAIN_SIG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN RIIO_BOND80x100_PLAIN_SIG 0 0 ;
  SIZE 80 BY 100 ;
  SYMMETRY X Y R90 ;
  SITE IO_BOND_site ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT 0 0 80 100 ;
    END
  END PAD
  OBS
    LAYER CA ;
      RECT 0 0 80 100 ;
    LAYER M1 ;
      RECT 0 0 80 100 ;
    LAYER V1 ;
      RECT 0 0 80 100 ;
    LAYER M2 ;
      RECT 0 0 80 100 ;
    LAYER A1 ;
      RECT 0 0 80 100 ;
    LAYER C2 ;
      RECT 0 0 80 100 ;
    LAYER IA ;
      RECT 0 0 80 100 ;
    LAYER LB ;
      RECT 0 0 80 100 ;
    LAYER VV ;
      RECT 0 0 80 100 ;
    LAYER XA ;
      RECT 0 0 80 100 ;
    LAYER YX ;
      RECT 0 0 80 100 ;
    LAYER IB ;
      RECT 0 0 80 100 ;
    LAYER CB ;
      RECT 0 0 80 100 ;
    LAYER AY ;
      RECT 0 0 80 100 ;
    LAYER C1 ;
      RECT 0 0 80 100 ;
    LAYER C5 ;
      RECT 0 0 80 100 ;
    LAYER C4 ;
      RECT 0 0 80 100 ;
    LAYER C3 ;
      RECT 0 0 80 100 ;
    LAYER A5 ;
      RECT 0 0 80 100 ;
    LAYER A4 ;
      RECT 0 0 80 100 ;
    LAYER A3 ;
      RECT 0 0 80 100 ;
    LAYER A2 ;
      RECT 0 0 80 100 ;
    LAYER C6 ;
      RECT 0 0 80 100 ;
  END
END RIIO_BOND80x100_PLAIN_SIG

MACRO RIIO_BUMP_RCUP100_DY
  CLASS COVER BUMP ;
  ORIGIN 30 30 ;
  FOREIGN RIIO_BUMP_RCUP100_DY -30 -30 ;
  SIZE 60.000 BY 60.000 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT -12.426 -30 12.426 30 ;
        RECT -30 -12.426 30 12.426 ;
    END
  END PAD
  OBS
    LAYER LB ;
      RECT -30.000 -14.183 30.000 14.183 ;
      RECT -28.243 -15.941 28.243 15.941 ;
      RECT -26.485 -17.698 26.485 17.698 ;
      RECT -24.728 -19.456 24.728 19.456 ;
      RECT -22.970 -21.213 22.970 21.213 ;
      RECT -21.213 -22.970 21.213 22.970 ;
      RECT -19.456 -24.728 19.456 24.728 ;
      RECT -17.698 -26.485 17.698 26.485 ;
      RECT -15.941 -28.243 15.941 28.243 ;
      RECT -14.183 -30.000 14.183 30.000 ;
    LAYER VV ;
      RECT -30.000 -14.183 30.000 14.183 ;
      RECT -28.243 -15.941 28.243 15.941 ;
      RECT -26.485 -17.698 26.485 17.698 ;
      RECT -24.728 -19.456 24.728 19.456 ;
      RECT -22.970 -21.213 22.970 21.213 ;
      RECT -21.213 -22.970 21.213 22.970 ;
      RECT -19.456 -24.728 19.456 24.728 ;
      RECT -17.698 -26.485 17.698 26.485 ;
      RECT -15.941 -28.243 15.941 28.243 ;
      RECT -14.183 -30.000 14.183 30.000 ;
  END
END RIIO_BUMP_RCUP100_DY
MACRO RIIO_BUMP_RCUP100_GND
  CLASS COVER BUMP ;
  ORIGIN 30 30 ;
  FOREIGN RIIO_BUMP_RCUP100_GND -30 -30 ;
  SIZE 60.000 BY 60.000 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
      RECT -30.000 -12.426 -1.030 12.426 ;
      RECT 1.030 -12.426 30.000 12.426 ;
      RECT -30.000 -12.426 30.000 -11.030 ;
      RECT -28.243 -14.183 28.243 -11.030 ;
      RECT -26.485 -15.941 26.485 -11.030 ;
      RECT -24.728 -17.698 24.728 -11.030 ;
      RECT -22.970 -19.456 22.970 -11.030 ;
      RECT -21.213 -21.213 21.213 -11.030 ;
      RECT -19.456 -22.970 19.456 -11.030 ;
      RECT -17.698 -24.728 17.698 -11.030 ;
      RECT -15.941 -26.485 15.941 -11.030 ;
      RECT -14.183 -28.243 14.183 -11.030 ;
      RECT -12.426 -30.000 12.426 -11.030 ;
      RECT -30.000 -8.970 30.000 12.426 ;
      RECT -28.243 -8.970 28.243 14.183 ;
      RECT -26.485 -8.970 26.485 15.941 ;
      RECT -24.728 -8.970 24.728 17.698 ;
      RECT -22.970 -8.970 22.970 19.456 ;
      RECT -21.213 -8.970 21.213 21.213 ;
      RECT -19.456 -8.970 19.456 22.970 ;
      RECT -17.698 -8.970 17.698 24.728 ;
      RECT -15.941 -8.970 15.941 26.485 ;
      RECT -14.183 -8.970 14.183 28.243 ;
      RECT -12.426 -8.970 12.426 30.000 ;
    END
  END VSS
  OBS
    LAYER VV ;
      RECT -30.000 -14.183 30.000 14.183 ;
      RECT -28.243 -15.941 28.243 15.941 ;
      RECT -26.485 -17.698 26.485 17.698 ;
      RECT -24.728 -19.456 24.728 19.456 ;
      RECT -22.970 -21.213 22.970 21.213 ;
      RECT -21.213 -22.970 21.213 22.970 ;
      RECT -19.456 -24.728 19.456 24.728 ;
      RECT -17.698 -26.485 17.698 26.485 ;
      RECT -15.941 -28.243 15.941 28.243 ;
      RECT -14.183 -30.000 14.183 30.000 ;
  END
END RIIO_BUMP_RCUP100_GND
MACRO RIIO_BUMP_RCUP100_PWR
  CLASS COVER BUMP ;
  ORIGIN 30 30 ;
  FOREIGN RIIO_BUMP_RCUP100_PWR -30 -30 ;
  SIZE 60.000 BY 60.000 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
      RECT -30.000 -12.426 -1.030 12.426 ;
      RECT 1.030 -12.426 30.000 12.426 ;
      RECT -30.000 -12.426 30.000 -11.030 ;
      RECT -28.243 -14.183 28.243 -11.030 ;
      RECT -26.485 -15.941 26.485 -11.030 ;
      RECT -24.728 -17.698 24.728 -11.030 ;
      RECT -22.970 -19.456 22.970 -11.030 ;
      RECT -21.213 -21.213 21.213 -11.030 ;
      RECT -19.456 -22.970 19.456 -11.030 ;
      RECT -17.698 -24.728 17.698 -11.030 ;
      RECT -15.941 -26.485 15.941 -11.030 ;
      RECT -14.183 -28.243 14.183 -11.030 ;
      RECT -12.426 -30.000 12.426 -11.030 ;
      RECT -30.000 -8.970 30.000 12.426 ;
      RECT -28.243 -8.970 28.243 14.183 ;
      RECT -26.485 -8.970 26.485 15.941 ;
      RECT -24.728 -8.970 24.728 17.698 ;
      RECT -22.970 -8.970 22.970 19.456 ;
      RECT -21.213 -8.970 21.213 21.213 ;
      RECT -19.456 -8.970 19.456 22.970 ;
      RECT -17.698 -8.970 17.698 24.728 ;
      RECT -15.941 -8.970 15.941 26.485 ;
      RECT -14.183 -8.970 14.183 28.243 ;
      RECT -12.426 -8.970 12.426 30.000 ;
    END
  END VDD
  OBS
    LAYER VV ;
      RECT -30.000 -14.183 30.000 14.183 ;
      RECT -28.243 -15.941 28.243 15.941 ;
      RECT -26.485 -17.698 26.485 17.698 ;
      RECT -24.728 -19.456 24.728 19.456 ;
      RECT -22.970 -21.213 22.970 21.213 ;
      RECT -21.213 -22.970 21.213 22.970 ;
      RECT -19.456 -24.728 19.456 24.728 ;
      RECT -17.698 -26.485 17.698 26.485 ;
      RECT -15.941 -28.243 15.941 28.243 ;
      RECT -14.183 -30.000 14.183 30.000 ;
  END
END RIIO_BUMP_RCUP100_PWR
MACRO RIIO_BUMP_RCUP100_SIG
  CLASS COVER BUMP ;
  ORIGIN 30 30 ;
  FOREIGN RIIO_BUMP_RCUP100_SIG -30 -30 ;
  SIZE 60.000 BY 60.000 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
      RECT -30.000 -12.426 -1.030 12.426 ;
      RECT 1.030 -12.426 30.000 12.426 ;
      RECT -30.000 -12.426 30.000 -11.030 ;
      RECT -28.243 -14.183 28.243 -11.030 ;
      RECT -26.485 -15.941 26.485 -11.030 ;
      RECT -24.728 -17.698 24.728 -11.030 ;
      RECT -22.970 -19.456 22.970 -11.030 ;
      RECT -21.213 -21.213 21.213 -11.030 ;
      RECT -19.456 -22.970 19.456 -11.030 ;
      RECT -17.698 -24.728 17.698 -11.030 ;
      RECT -15.941 -26.485 15.941 -11.030 ;
      RECT -14.183 -28.243 14.183 -11.030 ;
      RECT -12.426 -30.000 12.426 -11.030 ;
      RECT -30.000 -8.970 30.000 12.426 ;
      RECT -28.243 -8.970 28.243 14.183 ;
      RECT -26.485 -8.970 26.485 15.941 ;
      RECT -24.728 -8.970 24.728 17.698 ;
      RECT -22.970 -8.970 22.970 19.456 ;
      RECT -21.213 -8.970 21.213 21.213 ;
      RECT -19.456 -8.970 19.456 22.970 ;
      RECT -17.698 -8.970 17.698 24.728 ;
      RECT -15.941 -8.970 15.941 26.485 ;
      RECT -14.183 -8.970 14.183 28.243 ;
      RECT -12.426 -8.970 12.426 30.000 ;
    END
  END PAD
  OBS
    LAYER VV ;
      RECT -30.000 -14.183 30.000 14.183 ;
      RECT -28.243 -15.941 28.243 15.941 ;
      RECT -26.485 -17.698 26.485 17.698 ;
      RECT -24.728 -19.456 24.728 19.456 ;
      RECT -22.970 -21.213 22.970 21.213 ;
      RECT -21.213 -22.970 21.213 22.970 ;
      RECT -19.456 -24.728 19.456 24.728 ;
      RECT -17.698 -26.485 17.698 26.485 ;
      RECT -15.941 -28.243 15.941 28.243 ;
      RECT -14.183 -30.000 14.183 30.000 ;
  END
END RIIO_BUMP_RCUP100_SIG
MACRO RIIO_BUMP_RCUP130_DY
  CLASS COVER BUMP ;
  ORIGIN 45 45 ;
  FOREIGN RIIO_BUMP_RCUP130_DY -45 -45 ;
  SIZE 90.000 BY 90.000 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT -18.639 -45 18.639 45 ;
        RECT -45 -18.639 45 18.639 ;
    END
  END PAD
  OBS
    LAYER LB ;
      RECT -45.000 -21.275 45.000 21.275 ;
      RECT -42.364 -23.911 42.364 23.911 ;
      RECT -39.728 -26.547 39.728 26.547 ;
      RECT -37.092 -29.183 37.092 29.183 ;
      RECT -34.456 -31.820 34.456 31.820 ;
      RECT -31.819 -34.456 31.819 34.456 ;
      RECT -29.183 -37.092 29.183 37.092 ;
      RECT -26.547 -39.728 26.547 39.728 ;
      RECT -23.911 -42.364 23.911 42.364 ;
      RECT -21.275 -45.000 21.275 45.000 ;
    LAYER VV ;
      RECT -45.000 -21.275 45.000 21.275 ;
      RECT -42.364 -23.911 42.364 23.911 ;
      RECT -39.728 -26.547 39.728 26.547 ;
      RECT -37.092 -29.183 37.092 29.183 ;
      RECT -34.456 -31.820 34.456 31.820 ;
      RECT -31.819 -34.456 31.819 34.456 ;
      RECT -29.183 -37.092 29.183 37.092 ;
      RECT -26.547 -39.728 26.547 39.728 ;
      RECT -23.911 -42.364 23.911 42.364 ;
      RECT -21.275 -45.000 21.275 45.000 ;
  END
END RIIO_BUMP_RCUP130_DY
MACRO RIIO_BUMP_RCUP130_GND
  CLASS COVER BUMP ;
  ORIGIN 45 45 ;
  FOREIGN RIIO_BUMP_RCUP130_GND -45 -45 ;
  SIZE 90.000 BY 90.000 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
      RECT -45.000 -18.639 -1.030 18.639 ;
      RECT 1.030 -18.639 45.000 18.639 ;
      RECT -45.000 -18.639 45.000 -11.030 ;
      RECT -42.364 -21.275 42.364 -11.030 ;
      RECT -39.728 -23.911 39.728 -11.030 ;
      RECT -37.092 -26.547 37.092 -11.030 ;
      RECT -34.456 -29.183 34.456 -11.030 ;
      RECT -31.819 -31.820 31.819 -11.030 ;
      RECT -29.183 -34.456 29.183 -11.030 ;
      RECT -26.547 -37.092 26.547 -11.030 ;
      RECT -23.911 -39.728 23.911 -11.030 ;
      RECT -21.275 -42.364 21.275 -11.030 ;
      RECT -18.639 -45.000 18.639 -11.030 ;
      RECT -45.000 -8.970 45.000 18.639 ;
      RECT -42.364 -8.970 42.364 21.275 ;
      RECT -39.728 -8.970 39.728 23.911 ;
      RECT -37.092 -8.970 37.092 26.547 ;
      RECT -34.456 -8.970 34.456 29.183 ;
      RECT -31.819 -8.970 31.819 31.820 ;
      RECT -29.183 -8.970 29.183 34.456 ;
      RECT -26.547 -8.970 26.547 37.092 ;
      RECT -23.911 -8.970 23.911 39.728 ;
      RECT -21.275 -8.970 21.275 42.364 ;
      RECT -18.639 -8.970 18.639 45.000 ;
    END
  END VSS
  OBS
    LAYER VV ;
      RECT -45.000 -21.275 45.000 21.275 ;
      RECT -42.364 -23.911 42.364 23.911 ;
      RECT -39.728 -26.547 39.728 26.547 ;
      RECT -37.092 -29.183 37.092 29.183 ;
      RECT -34.456 -31.820 34.456 31.820 ;
      RECT -31.819 -34.456 31.819 34.456 ;
      RECT -29.183 -37.092 29.183 37.092 ;
      RECT -26.547 -39.728 26.547 39.728 ;
      RECT -23.911 -42.364 23.911 42.364 ;
      RECT -21.275 -45.000 21.275 45.000 ;
  END
END RIIO_BUMP_RCUP130_GND
MACRO RIIO_BUMP_RCUP130_PWR
  CLASS COVER BUMP ;
  ORIGIN 45 45 ;
  FOREIGN RIIO_BUMP_RCUP130_PWR -45 -45 ;
  SIZE 90.000 BY 90.000 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
      RECT -45.000 -18.639 -1.030 18.639 ;
      RECT 1.030 -18.639 45.000 18.639 ;
      RECT -45.000 -18.639 45.000 -11.030 ;
      RECT -42.364 -21.275 42.364 -11.030 ;
      RECT -39.728 -23.911 39.728 -11.030 ;
      RECT -37.092 -26.547 37.092 -11.030 ;
      RECT -34.456 -29.183 34.456 -11.030 ;
      RECT -31.819 -31.820 31.819 -11.030 ;
      RECT -29.183 -34.456 29.183 -11.030 ;
      RECT -26.547 -37.092 26.547 -11.030 ;
      RECT -23.911 -39.728 23.911 -11.030 ;
      RECT -21.275 -42.364 21.275 -11.030 ;
      RECT -18.639 -45.000 18.639 -11.030 ;
      RECT -45.000 -8.970 45.000 18.639 ;
      RECT -42.364 -8.970 42.364 21.275 ;
      RECT -39.728 -8.970 39.728 23.911 ;
      RECT -37.092 -8.970 37.092 26.547 ;
      RECT -34.456 -8.970 34.456 29.183 ;
      RECT -31.819 -8.970 31.819 31.820 ;
      RECT -29.183 -8.970 29.183 34.456 ;
      RECT -26.547 -8.970 26.547 37.092 ;
      RECT -23.911 -8.970 23.911 39.728 ;
      RECT -21.275 -8.970 21.275 42.364 ;
      RECT -18.639 -8.970 18.639 45.000 ;
    END
  END VDD
  OBS
    LAYER VV ;
      RECT -45.000 -21.275 45.000 21.275 ;
      RECT -42.364 -23.911 42.364 23.911 ;
      RECT -39.728 -26.547 39.728 26.547 ;
      RECT -37.092 -29.183 37.092 29.183 ;
      RECT -34.456 -31.820 34.456 31.820 ;
      RECT -31.819 -34.456 31.819 34.456 ;
      RECT -29.183 -37.092 29.183 37.092 ;
      RECT -26.547 -39.728 26.547 39.728 ;
      RECT -23.911 -42.364 23.911 42.364 ;
      RECT -21.275 -45.000 21.275 45.000 ;
  END
END RIIO_BUMP_RCUP130_PWR
MACRO RIIO_BUMP_RCUP130_SIG
  CLASS COVER BUMP ;
  ORIGIN 45 45 ;
  FOREIGN RIIO_BUMP_RCUP130_SIG -45 -45 ;
  SIZE 90.000 BY 90.000 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
      RECT -45.000 -18.639 -1.030 18.639 ;
      RECT 1.030 -18.639 45.000 18.639 ;
      RECT -45.000 -18.639 45.000 -11.030 ;
      RECT -42.364 -21.275 42.364 -11.030 ;
      RECT -39.728 -23.911 39.728 -11.030 ;
      RECT -37.092 -26.547 37.092 -11.030 ;
      RECT -34.456 -29.183 34.456 -11.030 ;
      RECT -31.819 -31.820 31.819 -11.030 ;
      RECT -29.183 -34.456 29.183 -11.030 ;
      RECT -26.547 -37.092 26.547 -11.030 ;
      RECT -23.911 -39.728 23.911 -11.030 ;
      RECT -21.275 -42.364 21.275 -11.030 ;
      RECT -18.639 -45.000 18.639 -11.030 ;
      RECT -45.000 -8.970 45.000 18.639 ;
      RECT -42.364 -8.970 42.364 21.275 ;
      RECT -39.728 -8.970 39.728 23.911 ;
      RECT -37.092 -8.970 37.092 26.547 ;
      RECT -34.456 -8.970 34.456 29.183 ;
      RECT -31.819 -8.970 31.819 31.820 ;
      RECT -29.183 -8.970 29.183 34.456 ;
      RECT -26.547 -8.970 26.547 37.092 ;
      RECT -23.911 -8.970 23.911 39.728 ;
      RECT -21.275 -8.970 21.275 42.364 ;
      RECT -18.639 -8.970 18.639 45.000 ;
    END
  END PAD
  OBS
    LAYER VV ;
      RECT -45.000 -21.275 45.000 21.275 ;
      RECT -42.364 -23.911 42.364 23.911 ;
      RECT -39.728 -26.547 39.728 26.547 ;
      RECT -37.092 -29.183 37.092 29.183 ;
      RECT -34.456 -31.820 34.456 31.820 ;
      RECT -31.819 -34.456 31.819 34.456 ;
      RECT -29.183 -37.092 29.183 37.092 ;
      RECT -26.547 -39.728 26.547 39.728 ;
      RECT -23.911 -42.364 23.911 42.364 ;
      RECT -21.275 -45.000 21.275 45.000 ;
  END
END RIIO_BUMP_RCUP130_SIG
MACRO RIIO_BUMP_SNAG140_DY
  CLASS COVER BUMP ;
  ORIGIN 35.5 35.5 ;
  FOREIGN RIIO_BUMP_SNAG140_DY -35.5 -35.5 ;
  SIZE 71.000 BY 71.000 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT -14.705 -35.5 14.705 35.5 ;
        RECT -35.5 -14.705 35.5 14.705 ;
    END
  END PAD
  OBS
    LAYER LB ;
      RECT -35.500 -16.784 35.500 16.784 ;
      RECT -33.420 -18.864 33.420 18.864 ;
      RECT -31.341 -20.944 31.341 20.944 ;
      RECT -29.261 -23.023 29.261 23.023 ;
      RECT -27.182 -25.102 27.182 25.102 ;
      RECT -25.103 -27.182 25.103 27.182 ;
      RECT -23.023 -29.261 23.023 29.261 ;
      RECT -20.944 -31.341 20.944 31.341 ;
      RECT -18.864 -33.420 18.864 33.420 ;
      RECT -16.785 -35.500 16.785 35.500 ;
    LAYER VV ;
      RECT -35.500 -16.784 35.500 16.784 ;
      RECT -33.420 -18.864 33.420 18.864 ;
      RECT -31.341 -20.944 31.341 20.944 ;
      RECT -29.261 -23.023 29.261 23.023 ;
      RECT -27.182 -25.102 27.182 25.102 ;
      RECT -25.103 -27.182 25.103 27.182 ;
      RECT -23.023 -29.261 23.023 29.261 ;
      RECT -20.944 -31.341 20.944 31.341 ;
      RECT -18.864 -33.420 18.864 33.420 ;
      RECT -16.785 -35.500 16.785 35.500 ;
  END
END RIIO_BUMP_SNAG140_DY
MACRO RIIO_BUMP_SNAG140_GND
  CLASS COVER BUMP ;
  ORIGIN 35.5 35.5 ;
  FOREIGN RIIO_BUMP_SNAG140_GND -35.5 -35.5 ;
  SIZE 71.000 BY 71.000 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
      RECT -35.500 -14.705 -1.030 14.705 ;
      RECT 1.030 -14.705 35.500 14.705 ;
      RECT -35.500 -14.705 35.500 -11.030 ;
      RECT -33.420 -16.784 33.420 -11.030 ;
      RECT -31.341 -18.864 31.341 -11.030 ;
      RECT -29.261 -20.944 29.261 -11.030 ;
      RECT -27.182 -23.023 27.182 -11.030 ;
      RECT -25.103 -25.102 25.103 -11.030 ;
      RECT -23.023 -27.182 23.023 -11.030 ;
      RECT -20.944 -29.261 20.944 -11.030 ;
      RECT -18.864 -31.341 18.864 -11.030 ;
      RECT -16.785 -33.420 16.785 -11.030 ;
      RECT -14.705 -35.500 14.705 -11.030 ;
      RECT -35.500 -8.970 35.500 14.705 ;
      RECT -33.420 -8.970 33.420 16.784 ;
      RECT -31.341 -8.970 31.341 18.864 ;
      RECT -29.261 -8.970 29.261 20.944 ;
      RECT -27.182 -8.970 27.182 23.023 ;
      RECT -25.103 -8.970 25.103 25.102 ;
      RECT -23.023 -8.970 23.023 27.182 ;
      RECT -20.944 -8.970 20.944 29.261 ;
      RECT -18.864 -8.970 18.864 31.341 ;
      RECT -16.785 -8.970 16.785 33.420 ;
      RECT -14.705 -8.970 14.705 35.500 ;
    END
  END VSS
  OBS
    LAYER VV ;
      RECT -35.500 -16.784 35.500 16.784 ;
      RECT -33.420 -18.864 33.420 18.864 ;
      RECT -31.341 -20.944 31.341 20.944 ;
      RECT -29.261 -23.023 29.261 23.023 ;
      RECT -27.182 -25.102 27.182 25.102 ;
      RECT -25.103 -27.182 25.103 27.182 ;
      RECT -23.023 -29.261 23.023 29.261 ;
      RECT -20.944 -31.341 20.944 31.341 ;
      RECT -18.864 -33.420 18.864 33.420 ;
      RECT -16.785 -35.500 16.785 35.500 ;
  END
END RIIO_BUMP_SNAG140_GND
MACRO RIIO_BUMP_SNAG140_PWR
  CLASS COVER BUMP ;
  ORIGIN 35.5 35.5 ;
  FOREIGN RIIO_BUMP_SNAG140_PWR -35.5 -35.5 ;
  SIZE 71.000 BY 71.000 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
      RECT -35.500 -14.705 -1.030 14.705 ;
      RECT 1.030 -14.705 35.500 14.705 ;
      RECT -35.500 -14.705 35.500 -11.030 ;
      RECT -33.420 -16.784 33.420 -11.030 ;
      RECT -31.341 -18.864 31.341 -11.030 ;
      RECT -29.261 -20.944 29.261 -11.030 ;
      RECT -27.182 -23.023 27.182 -11.030 ;
      RECT -25.103 -25.102 25.103 -11.030 ;
      RECT -23.023 -27.182 23.023 -11.030 ;
      RECT -20.944 -29.261 20.944 -11.030 ;
      RECT -18.864 -31.341 18.864 -11.030 ;
      RECT -16.785 -33.420 16.785 -11.030 ;
      RECT -14.705 -35.500 14.705 -11.030 ;
      RECT -35.500 -8.970 35.500 14.705 ;
      RECT -33.420 -8.970 33.420 16.784 ;
      RECT -31.341 -8.970 31.341 18.864 ;
      RECT -29.261 -8.970 29.261 20.944 ;
      RECT -27.182 -8.970 27.182 23.023 ;
      RECT -25.103 -8.970 25.103 25.102 ;
      RECT -23.023 -8.970 23.023 27.182 ;
      RECT -20.944 -8.970 20.944 29.261 ;
      RECT -18.864 -8.970 18.864 31.341 ;
      RECT -16.785 -8.970 16.785 33.420 ;
      RECT -14.705 -8.970 14.705 35.500 ;
    END
  END VDD
  OBS
    LAYER VV ;
      RECT -35.500 -16.784 35.500 16.784 ;
      RECT -33.420 -18.864 33.420 18.864 ;
      RECT -31.341 -20.944 31.341 20.944 ;
      RECT -29.261 -23.023 29.261 23.023 ;
      RECT -27.182 -25.102 27.182 25.102 ;
      RECT -25.103 -27.182 25.103 27.182 ;
      RECT -23.023 -29.261 23.023 29.261 ;
      RECT -20.944 -31.341 20.944 31.341 ;
      RECT -18.864 -33.420 18.864 33.420 ;
      RECT -16.785 -35.500 16.785 35.500 ;
  END
END RIIO_BUMP_SNAG140_PWR
MACRO RIIO_BUMP_SNAG140_SIG
  CLASS COVER BUMP ;
  ORIGIN 35.5 35.5 ;
  FOREIGN RIIO_BUMP_SNAG140_SIG -35.5 -35.5 ;
  SIZE 71.000 BY 71.000 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
      RECT -35.500 -14.705 -1.030 14.705 ;
      RECT 1.030 -14.705 35.500 14.705 ;
      RECT -35.500 -14.705 35.500 -11.030 ;
      RECT -33.420 -16.784 33.420 -11.030 ;
      RECT -31.341 -18.864 31.341 -11.030 ;
      RECT -29.261 -20.944 29.261 -11.030 ;
      RECT -27.182 -23.023 27.182 -11.030 ;
      RECT -25.103 -25.102 25.103 -11.030 ;
      RECT -23.023 -27.182 23.023 -11.030 ;
      RECT -20.944 -29.261 20.944 -11.030 ;
      RECT -18.864 -31.341 18.864 -11.030 ;
      RECT -16.785 -33.420 16.785 -11.030 ;
      RECT -14.705 -35.500 14.705 -11.030 ;
      RECT -35.500 -8.970 35.500 14.705 ;
      RECT -33.420 -8.970 33.420 16.784 ;
      RECT -31.341 -8.970 31.341 18.864 ;
      RECT -29.261 -8.970 29.261 20.944 ;
      RECT -27.182 -8.970 27.182 23.023 ;
      RECT -25.103 -8.970 25.103 25.102 ;
      RECT -23.023 -8.970 23.023 27.182 ;
      RECT -20.944 -8.970 20.944 29.261 ;
      RECT -18.864 -8.970 18.864 31.341 ;
      RECT -16.785 -8.970 16.785 33.420 ;
      RECT -14.705 -8.970 14.705 35.500 ;
    END
  END PAD
  OBS
    LAYER VV ;
      RECT -35.500 -16.784 35.500 16.784 ;
      RECT -33.420 -18.864 33.420 18.864 ;
      RECT -31.341 -20.944 31.341 20.944 ;
      RECT -29.261 -23.023 29.261 23.023 ;
      RECT -27.182 -25.102 27.182 25.102 ;
      RECT -25.103 -27.182 25.103 27.182 ;
      RECT -23.023 -29.261 23.023 29.261 ;
      RECT -20.944 -31.341 20.944 31.341 ;
      RECT -18.864 -33.420 18.864 33.420 ;
      RECT -16.785 -35.500 16.785 35.500 ;
  END
END RIIO_BUMP_SNAG140_SIG
MACRO RIIO_BUMP_SNAG150_DY
  CLASS COVER BUMP ;
  ORIGIN 40.8 40.8 ;
  FOREIGN RIIO_BUMP_SNAG150_DY -40.8 -40.8 ;
  SIZE 81.600 BY 81.600 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT -16.9 -40.8 16.9 40.8 ;
        RECT -40.8 -16.9 40.8 16.9 ;
    END
  END PAD
  OBS
    LAYER LB ;
      RECT -40.800 -19.290 40.800 19.290 ;
      RECT -38.410 -21.680 38.410 21.680 ;
      RECT -36.020 -24.070 36.020 24.070 ;
      RECT -33.630 -26.460 33.630 26.460 ;
      RECT -31.240 -28.850 31.240 28.850 ;
      RECT -28.850 -31.240 28.850 31.240 ;
      RECT -26.460 -33.630 26.460 33.630 ;
      RECT -24.070 -36.020 24.070 36.020 ;
      RECT -21.680 -38.410 21.680 38.410 ;
      RECT -19.290 -40.800 19.290 40.800 ;
    LAYER VV ;
      RECT -40.800 -19.290 40.800 19.290 ;
      RECT -38.410 -21.680 38.410 21.680 ;
      RECT -36.020 -24.070 36.020 24.070 ;
      RECT -33.630 -26.460 33.630 26.460 ;
      RECT -31.240 -28.850 31.240 28.850 ;
      RECT -28.850 -31.240 28.850 31.240 ;
      RECT -26.460 -33.630 26.460 33.630 ;
      RECT -24.070 -36.020 24.070 36.020 ;
      RECT -21.680 -38.410 21.680 38.410 ;
      RECT -19.290 -40.800 19.290 40.800 ;
  END
END RIIO_BUMP_SNAG150_DY
MACRO RIIO_BUMP_SNAG150_GND
  CLASS COVER BUMP ;
  ORIGIN 40.8 40.8 ;
  FOREIGN RIIO_BUMP_SNAG150_GND -40.8 -40.8 ;
  SIZE 81.600 BY 81.600 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
      RECT -40.800 -16.900 -1.030 16.900 ;
      RECT 1.030 -16.900 40.800 16.900 ;
      RECT -40.800 -16.900 40.800 -11.030 ;
      RECT -38.410 -19.290 38.410 -11.030 ;
      RECT -36.020 -21.680 36.020 -11.030 ;
      RECT -33.630 -24.070 33.630 -11.030 ;
      RECT -31.240 -26.460 31.240 -11.030 ;
      RECT -28.850 -28.850 28.850 -11.030 ;
      RECT -26.460 -31.240 26.460 -11.030 ;
      RECT -24.070 -33.630 24.070 -11.030 ;
      RECT -21.680 -36.020 21.680 -11.030 ;
      RECT -19.290 -38.410 19.290 -11.030 ;
      RECT -16.900 -40.800 16.900 -11.030 ;
      RECT -40.800 -8.970 40.800 16.900 ;
      RECT -38.410 -8.970 38.410 19.290 ;
      RECT -36.020 -8.970 36.020 21.680 ;
      RECT -33.630 -8.970 33.630 24.070 ;
      RECT -31.240 -8.970 31.240 26.460 ;
      RECT -28.850 -8.970 28.850 28.850 ;
      RECT -26.460 -8.970 26.460 31.240 ;
      RECT -24.070 -8.970 24.070 33.630 ;
      RECT -21.680 -8.970 21.680 36.020 ;
      RECT -19.290 -8.970 19.290 38.410 ;
      RECT -16.900 -8.970 16.900 40.800 ;
    END
  END VSS
  OBS
    LAYER VV ;
      RECT -40.800 -19.290 40.800 19.290 ;
      RECT -38.410 -21.680 38.410 21.680 ;
      RECT -36.020 -24.070 36.020 24.070 ;
      RECT -33.630 -26.460 33.630 26.460 ;
      RECT -31.240 -28.850 31.240 28.850 ;
      RECT -28.850 -31.240 28.850 31.240 ;
      RECT -26.460 -33.630 26.460 33.630 ;
      RECT -24.070 -36.020 24.070 36.020 ;
      RECT -21.680 -38.410 21.680 38.410 ;
      RECT -19.290 -40.800 19.290 40.800 ;
  END
END RIIO_BUMP_SNAG150_GND
MACRO RIIO_BUMP_SNAG150_PWR
  CLASS COVER BUMP ;
  ORIGIN 40.8 40.8 ;
  FOREIGN RIIO_BUMP_SNAG150_PWR -40.8 -40.8 ;
  SIZE 81.600 BY 81.600 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
      RECT -40.800 -16.900 -1.030 16.900 ;
      RECT 1.030 -16.900 40.800 16.900 ;
      RECT -40.800 -16.900 40.800 -11.030 ;
      RECT -38.410 -19.290 38.410 -11.030 ;
      RECT -36.020 -21.680 36.020 -11.030 ;
      RECT -33.630 -24.070 33.630 -11.030 ;
      RECT -31.240 -26.460 31.240 -11.030 ;
      RECT -28.850 -28.850 28.850 -11.030 ;
      RECT -26.460 -31.240 26.460 -11.030 ;
      RECT -24.070 -33.630 24.070 -11.030 ;
      RECT -21.680 -36.020 21.680 -11.030 ;
      RECT -19.290 -38.410 19.290 -11.030 ;
      RECT -16.900 -40.800 16.900 -11.030 ;
      RECT -40.800 -8.970 40.800 16.900 ;
      RECT -38.410 -8.970 38.410 19.290 ;
      RECT -36.020 -8.970 36.020 21.680 ;
      RECT -33.630 -8.970 33.630 24.070 ;
      RECT -31.240 -8.970 31.240 26.460 ;
      RECT -28.850 -8.970 28.850 28.850 ;
      RECT -26.460 -8.970 26.460 31.240 ;
      RECT -24.070 -8.970 24.070 33.630 ;
      RECT -21.680 -8.970 21.680 36.020 ;
      RECT -19.290 -8.970 19.290 38.410 ;
      RECT -16.900 -8.970 16.900 40.800 ;
    END
  END VDD
  OBS
    LAYER VV ;
      RECT -40.800 -19.290 40.800 19.290 ;
      RECT -38.410 -21.680 38.410 21.680 ;
      RECT -36.020 -24.070 36.020 24.070 ;
      RECT -33.630 -26.460 33.630 26.460 ;
      RECT -31.240 -28.850 31.240 28.850 ;
      RECT -28.850 -31.240 28.850 31.240 ;
      RECT -26.460 -33.630 26.460 33.630 ;
      RECT -24.070 -36.020 24.070 36.020 ;
      RECT -21.680 -38.410 21.680 38.410 ;
      RECT -19.290 -40.800 19.290 40.800 ;
  END
END RIIO_BUMP_SNAG150_PWR
MACRO RIIO_BUMP_SNAG150_SIG
  CLASS COVER BUMP ;
  ORIGIN 40.8 40.8 ;
  FOREIGN RIIO_BUMP_SNAG150_SIG -40.8 -40.8 ;
  SIZE 81.600 BY 81.600 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
      RECT -40.800 -16.900 -1.030 16.900 ;
      RECT 1.030 -16.900 40.800 16.900 ;
      RECT -40.800 -16.900 40.800 -11.030 ;
      RECT -38.410 -19.290 38.410 -11.030 ;
      RECT -36.020 -21.680 36.020 -11.030 ;
      RECT -33.630 -24.070 33.630 -11.030 ;
      RECT -31.240 -26.460 31.240 -11.030 ;
      RECT -28.850 -28.850 28.850 -11.030 ;
      RECT -26.460 -31.240 26.460 -11.030 ;
      RECT -24.070 -33.630 24.070 -11.030 ;
      RECT -21.680 -36.020 21.680 -11.030 ;
      RECT -19.290 -38.410 19.290 -11.030 ;
      RECT -16.900 -40.800 16.900 -11.030 ;
      RECT -40.800 -8.970 40.800 16.900 ;
      RECT -38.410 -8.970 38.410 19.290 ;
      RECT -36.020 -8.970 36.020 21.680 ;
      RECT -33.630 -8.970 33.630 24.070 ;
      RECT -31.240 -8.970 31.240 26.460 ;
      RECT -28.850 -8.970 28.850 28.850 ;
      RECT -26.460 -8.970 26.460 31.240 ;
      RECT -24.070 -8.970 24.070 33.630 ;
      RECT -21.680 -8.970 21.680 36.020 ;
      RECT -19.290 -8.970 19.290 38.410 ;
      RECT -16.900 -8.970 16.900 40.800 ;
    END
  END PAD
  OBS
    LAYER VV ;
      RECT -40.800 -19.290 40.800 19.290 ;
      RECT -38.410 -21.680 38.410 21.680 ;
      RECT -36.020 -24.070 36.020 24.070 ;
      RECT -33.630 -26.460 33.630 26.460 ;
      RECT -31.240 -28.850 31.240 28.850 ;
      RECT -28.850 -31.240 28.850 31.240 ;
      RECT -26.460 -33.630 26.460 33.630 ;
      RECT -24.070 -36.020 24.070 36.020 ;
      RECT -21.680 -38.410 21.680 38.410 ;
      RECT -19.290 -40.800 19.290 40.800 ;
  END
END RIIO_BUMP_SNAG150_SIG
MACRO RIIO_BUMP_SNAG180_DY
  CLASS COVER BUMP ;
  ORIGIN 48 48 ;
  FOREIGN RIIO_BUMP_SNAG180_DY -48 -48 ;
  SIZE 96.000 BY 96.000 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
        RECT -19.882 -48 19.882 48 ;
        RECT -48 -19.882 48 19.882 ;
    END
  END PAD
  OBS
    LAYER LB ;
      RECT -48.000 -22.694 48.000 22.694 ;
      RECT -45.188 -25.506 45.188 25.506 ;
      RECT -42.376 -28.317 42.376 28.317 ;
      RECT -39.565 -31.129 39.565 31.129 ;
      RECT -36.753 -33.941 36.753 33.941 ;
      RECT -33.941 -36.753 33.941 36.753 ;
      RECT -31.129 -39.565 31.129 39.565 ;
      RECT -28.317 -42.376 28.317 42.376 ;
      RECT -25.506 -45.188 25.506 45.188 ;
      RECT -22.694 -48.000 22.694 48.000 ;
    LAYER VV ;
      RECT -48.000 -22.694 48.000 22.694 ;
      RECT -45.188 -25.506 45.188 25.506 ;
      RECT -42.376 -28.317 42.376 28.317 ;
      RECT -39.565 -31.129 39.565 31.129 ;
      RECT -36.753 -33.941 36.753 33.941 ;
      RECT -33.941 -36.753 33.941 36.753 ;
      RECT -31.129 -39.565 31.129 39.565 ;
      RECT -28.317 -42.376 28.317 42.376 ;
      RECT -25.506 -45.188 25.506 45.188 ;
      RECT -22.694 -48.000 22.694 48.000 ;
  END
END RIIO_BUMP_SNAG180_DY
MACRO RIIO_BUMP_SNAG180_GND
  CLASS COVER BUMP ;
  ORIGIN 48 48 ;
  FOREIGN RIIO_BUMP_SNAG180_GND -48 -48 ;
  SIZE 96.000 BY 96.000 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER LB ;
      RECT -48.000 -19.882 -1.030 19.882 ;
      RECT 1.030 -19.882 48.000 19.882 ;
      RECT -48.000 -19.882 48.000 -11.030 ;
      RECT -45.188 -22.694 45.188 -11.030 ;
      RECT -42.376 -25.506 42.376 -11.030 ;
      RECT -39.565 -28.317 39.565 -11.030 ;
      RECT -36.753 -31.129 36.753 -11.030 ;
      RECT -33.941 -33.941 33.941 -11.030 ;
      RECT -31.129 -36.753 31.129 -11.030 ;
      RECT -28.317 -39.565 28.317 -11.030 ;
      RECT -25.506 -42.376 25.506 -11.030 ;
      RECT -22.694 -45.188 22.694 -11.030 ;
      RECT -19.882 -48.000 19.882 -11.030 ;
      RECT -48.000 -8.970 48.000 19.882 ;
      RECT -45.188 -8.970 45.188 22.694 ;
      RECT -42.376 -8.970 42.376 25.506 ;
      RECT -39.565 -8.970 39.565 28.317 ;
      RECT -36.753 -8.970 36.753 31.129 ;
      RECT -33.941 -8.970 33.941 33.941 ;
      RECT -31.129 -8.970 31.129 36.753 ;
      RECT -28.317 -8.970 28.317 39.565 ;
      RECT -25.506 -8.970 25.506 42.376 ;
      RECT -22.694 -8.970 22.694 45.188 ;
      RECT -19.882 -8.970 19.882 48.000 ;
    END
  END VSS
  OBS
    LAYER VV ;
      RECT -48.000 -22.694 48.000 22.694 ;
      RECT -45.188 -25.506 45.188 25.506 ;
      RECT -42.376 -28.317 42.376 28.317 ;
      RECT -39.565 -31.129 39.565 31.129 ;
      RECT -36.753 -33.941 36.753 33.941 ;
      RECT -33.941 -36.753 33.941 36.753 ;
      RECT -31.129 -39.565 31.129 39.565 ;
      RECT -28.317 -42.376 28.317 42.376 ;
      RECT -25.506 -45.188 25.506 45.188 ;
      RECT -22.694 -48.000 22.694 48.000 ;
  END
END RIIO_BUMP_SNAG180_GND
MACRO RIIO_BUMP_SNAG180_PWR
  CLASS COVER BUMP ;
  ORIGIN 48 48 ;
  FOREIGN RIIO_BUMP_SNAG180_PWR -48 -48 ;
  SIZE 96.000 BY 96.000 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER LB ;
      RECT -48.000 -19.882 -1.030 19.882 ;
      RECT 1.030 -19.882 48.000 19.882 ;
      RECT -48.000 -19.882 48.000 -11.030 ;
      RECT -45.188 -22.694 45.188 -11.030 ;
      RECT -42.376 -25.506 42.376 -11.030 ;
      RECT -39.565 -28.317 39.565 -11.030 ;
      RECT -36.753 -31.129 36.753 -11.030 ;
      RECT -33.941 -33.941 33.941 -11.030 ;
      RECT -31.129 -36.753 31.129 -11.030 ;
      RECT -28.317 -39.565 28.317 -11.030 ;
      RECT -25.506 -42.376 25.506 -11.030 ;
      RECT -22.694 -45.188 22.694 -11.030 ;
      RECT -19.882 -48.000 19.882 -11.030 ;
      RECT -48.000 -8.970 48.000 19.882 ;
      RECT -45.188 -8.970 45.188 22.694 ;
      RECT -42.376 -8.970 42.376 25.506 ;
      RECT -39.565 -8.970 39.565 28.317 ;
      RECT -36.753 -8.970 36.753 31.129 ;
      RECT -33.941 -8.970 33.941 33.941 ;
      RECT -31.129 -8.970 31.129 36.753 ;
      RECT -28.317 -8.970 28.317 39.565 ;
      RECT -25.506 -8.970 25.506 42.376 ;
      RECT -22.694 -8.970 22.694 45.188 ;
      RECT -19.882 -8.970 19.882 48.000 ;
    END
  END VDD
  OBS
    LAYER VV ;
      RECT -48.000 -22.694 48.000 22.694 ;
      RECT -45.188 -25.506 45.188 25.506 ;
      RECT -42.376 -28.317 42.376 28.317 ;
      RECT -39.565 -31.129 39.565 31.129 ;
      RECT -36.753 -33.941 36.753 33.941 ;
      RECT -33.941 -36.753 33.941 36.753 ;
      RECT -31.129 -39.565 31.129 39.565 ;
      RECT -28.317 -42.376 28.317 42.376 ;
      RECT -25.506 -45.188 25.506 45.188 ;
      RECT -22.694 -48.000 22.694 48.000 ;
  END
END RIIO_BUMP_SNAG180_PWR
MACRO RIIO_BUMP_SNAG180_SIG
  CLASS COVER BUMP ;
  ORIGIN 48 48 ;
  FOREIGN RIIO_BUMP_SNAG180_SIG -48 -48 ;
  SIZE 96.000 BY 96.000 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER LB ;
      RECT -48.000 -19.882 -1.030 19.882 ;
      RECT 1.030 -19.882 48.000 19.882 ;
      RECT -48.000 -19.882 48.000 -11.030 ;
      RECT -45.188 -22.694 45.188 -11.030 ;
      RECT -42.376 -25.506 42.376 -11.030 ;
      RECT -39.565 -28.317 39.565 -11.030 ;
      RECT -36.753 -31.129 36.753 -11.030 ;
      RECT -33.941 -33.941 33.941 -11.030 ;
      RECT -31.129 -36.753 31.129 -11.030 ;
      RECT -28.317 -39.565 28.317 -11.030 ;
      RECT -25.506 -42.376 25.506 -11.030 ;
      RECT -22.694 -45.188 22.694 -11.030 ;
      RECT -19.882 -48.000 19.882 -11.030 ;
      RECT -48.000 -8.970 48.000 19.882 ;
      RECT -45.188 -8.970 45.188 22.694 ;
      RECT -42.376 -8.970 42.376 25.506 ;
      RECT -39.565 -8.970 39.565 28.317 ;
      RECT -36.753 -8.970 36.753 31.129 ;
      RECT -33.941 -8.970 33.941 33.941 ;
      RECT -31.129 -8.970 31.129 36.753 ;
      RECT -28.317 -8.970 28.317 39.565 ;
      RECT -25.506 -8.970 25.506 42.376 ;
      RECT -22.694 -8.970 22.694 45.188 ;
      RECT -19.882 -8.970 19.882 48.000 ;
    END
  END PAD
  OBS
    LAYER VV ;
      RECT -48.000 -22.694 48.000 22.694 ;
      RECT -45.188 -25.506 45.188 25.506 ;
      RECT -42.376 -28.317 42.376 28.317 ;
      RECT -39.565 -31.129 39.565 31.129 ;
      RECT -36.753 -33.941 36.753 33.941 ;
      RECT -33.941 -36.753 33.941 36.753 ;
      RECT -31.129 -39.565 31.129 39.565 ;
      RECT -28.317 -42.376 28.317 42.376 ;
      RECT -25.506 -45.188 25.506 45.188 ;
      RECT -22.694 -48.000 22.694 48.000 ;
  END
END RIIO_BUMP_SNAG180_SIG
END LIBRARY
